// Benchmark "c2670_blif" written by ABC on Sun Apr 14 20:10:46 2019

module c2670_blif  ( 
    G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
    G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
    G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
    G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
    G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
    G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
    G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136,
    G137, G138, G139, G140, G141, G142, ING169 , ING174 , ING177 ,
    ING178 , ING179 , ING180 , ING181 , ING182 , ING183 ,
    ING184 , ING185 , ING186 , ING189 , ING190 , ING191 ,
    ING192 , ING193 , ING194 , ING195 , ING196 , ING197 ,
    ING198 , ING199 , ING200 , ING201 , ING202 , ING203 ,
    ING204 , ING205 , ING206 , ING207 , ING208 , ING209 ,
    ING210 , ING211 , ING212 , ING213 , ING214 , ING215 ,
    ING239 , ING240 , ING241 , ING242 , ING243 , ING244 ,
    ING245 , ING246 , ING247 , ING248 , ING249 , ING250 ,
    ING251 , ING252 , ING253 , ING254 , ING255 , ING256 ,
    ING257 , ING262 , ING263 , ING264 , ING265 , ING266 ,
    ING267 , ING268 , ING269 , ING270 , ING271 , ING272 ,
    ING273 , ING274 , ING275 , ING276 , ING277 , ING278 ,
    ING279 , G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083,
    G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986,
    G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100,
    G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451,
    G2454, G2474, G2678,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G350, G335, G409, G369, G367, G411, G337, G384,
    G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173,
    G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171,
    G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
    G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145,
    G395, G295, G331, G397, G329, G231, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20,
    G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36,
    G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74,
    G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90,
    G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105,
    G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
    G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135,
    G136, G137, G138, G139, G140, G141, G142, ING169 , ING174 ,
    ING177 , ING178 , ING179 , ING180 , ING181 , ING182 ,
    ING183 , ING184 , ING185 , ING186 , ING189 , ING190 ,
    ING191 , ING192 , ING193 , ING194 , ING195 , ING196 ,
    ING197 , ING198 , ING199 , ING200 , ING201 , ING202 ,
    ING203 , ING204 , ING205 , ING206 , ING207 , ING208 ,
    ING209 , ING210 , ING211 , ING212 , ING213 , ING214 ,
    ING215 , ING239 , ING240 , ING241 , ING242 , ING243 ,
    ING244 , ING245 , ING246 , ING247 , ING248 , ING249 ,
    ING250 , ING251 , ING252 , ING253 , ING254 , ING255 ,
    ING256 , ING257 , ING262 , ING263 , ING264 , ING265 ,
    ING266 , ING267 , ING268 , ING269 , ING270 , ING271 ,
    ING272 , ING273 , ING274 , ING275 , ING276 , ING277 ,
    ING278 , ING279 , G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185,
    G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199,
    G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211,
    G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
    G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262,
    G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274,
    G275, G276, G277, G278, G279, G350, G335, G409, G369, G367, G411, G337,
    G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391,
    G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168,
    G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284,
    G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
    G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire n382, n383, n384, n385, n386, n387, n388, n389, n390, n392, n393,
    n394, n395, n396, n397, n399, n400, n402, n403, n405, n406, n408, n409,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n425, n426, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n446, n447, n448, n449, n450,
    n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n462, n463,
    n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
    n476, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523, n524, n525, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n546, n547, n548, n549, n550, n551, n552, n553, n555, n556,
    n557, n558, n559, n560, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n588, n589, n590, n591, n592, n593, n594, n595,
    n596, n597, n598, n599, n600, n601, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615, n616, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n637, n638, n640, n641, n642, n644, n645, n646, n647, n648,
    n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n673, n674,
    n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717, n718, n719, n721, n722, n723,
    n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
    n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791, n792, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
    n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
    n1043, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
    n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
    n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327;
  inv1   g0000(.a(G44), .O(G218));
  inv1   g0001(.a(G132), .O(G219));
  inv1   g0002(.a(G82), .O(G220));
  inv1   g0003(.a(G96), .O(G221));
  inv1   g0004(.a(G69), .O(G235));
  inv1   g0005(.a(G120), .O(G236));
  inv1   g0006(.a(G57), .O(G237));
  inv1   g0007(.a(G108), .O(G238));
  inv1   g0008(.a(G2072), .O(n382));
  inv1   g0009(.a(G2078), .O(n383));
  nor2   g0010(.a(n383), .b(n382), .O(n384));
  inv1   g0011(.a(n384), .O(n385));
  inv1   g0012(.a(G2084), .O(n386));
  inv1   g0013(.a(G2090), .O(n387));
  nor2   g0014(.a(n387), .b(n386), .O(n388));
  inv1   g0015(.a(n388), .O(n389));
  nor2   g0016(.a(n389), .b(n385), .O(n390));
  inv1   g0017(.a(n390), .O(G158));
  inv1   g0018(.a(G661), .O(n392));
  inv1   g0019(.a(G2), .O(n393));
  inv1   g0020(.a(G15), .O(n394));
  nor2   g0021(.a(n394), .b(n393), .O(n395));
  inv1   g0022(.a(n395), .O(n396));
  nor2   g0023(.a(n396), .b(n392), .O(n397));
  inv1   g0024(.a(n397), .O(G259));
  inv1   g0025(.a(G94), .O(n399));
  inv1   g0026(.a(G452), .O(n400));
  nor2   g0027(.a(n400), .b(n399), .O(G173));
  inv1   g0028(.a(G7), .O(n402));
  nor2   g0029(.a(n392), .b(n402), .O(n403));
  inv1   g0030(.a(n403), .O(G223));
  inv1   g0031(.a(G567), .O(n405));
  nor2   g0032(.a(G223), .b(n405), .O(n406));
  inv1   g0033(.a(n406), .O(G234));
  inv1   g0034(.a(G2106), .O(n408));
  nor2   g0035(.a(G223), .b(n408), .O(n409));
  inv1   g0036(.a(n409), .O(G217));
  nor2   g0037(.a(G235), .b(G237), .O(n411));
  inv1   g0038(.a(n411), .O(n412));
  nor2   g0039(.a(G236), .b(G238), .O(n413));
  inv1   g0040(.a(n413), .O(n414));
  nor2   g0041(.a(n414), .b(n412), .O(n415));
  inv1   g0042(.a(n415), .O(n416));
  nor2   g0043(.a(G220), .b(G218), .O(n417));
  inv1   g0044(.a(n417), .O(n418));
  nor2   g0045(.a(G219), .b(G221), .O(n419));
  inv1   g0046(.a(n419), .O(n420));
  nor2   g0047(.a(n420), .b(n418), .O(n421));
  inv1   g0048(.a(n421), .O(n422));
  nor2   g0049(.a(n422), .b(n416), .O(G325));
  inv1   g0050(.a(G325), .O(G261));
  nor2   g0051(.a(n421), .b(n408), .O(n425));
  nor2   g0052(.a(n415), .b(n405), .O(n426));
  nor2   g0053(.a(n426), .b(n425), .O(G319));
  inv1   g0054(.a(G113), .O(n428));
  inv1   g0055(.a(G2104), .O(n429));
  nor2   g0056(.a(n429), .b(n428), .O(n430));
  inv1   g0057(.a(G2105), .O(n431));
  inv1   g0058(.a(G125), .O(n432));
  nor2   g0059(.a(G2104), .b(n432), .O(n433));
  nor2   g0060(.a(n433), .b(n431), .O(n434));
  inv1   g0061(.a(n434), .O(n435));
  nor2   g0062(.a(n435), .b(n430), .O(n436));
  inv1   g0063(.a(G101), .O(n437));
  nor2   g0064(.a(n429), .b(n437), .O(n438));
  inv1   g0065(.a(G137), .O(n439));
  nor2   g0066(.a(G2104), .b(n439), .O(n440));
  nor2   g0067(.a(n440), .b(G2105), .O(n441));
  inv1   g0068(.a(n441), .O(n442));
  nor2   g0069(.a(n442), .b(n438), .O(n443));
  nor2   g0070(.a(n443), .b(n436), .O(n444));
  inv1   g0071(.a(n444), .O(G160));
  inv1   g0072(.a(G112), .O(n446));
  nor2   g0073(.a(n429), .b(n446), .O(n447));
  inv1   g0074(.a(G124), .O(n448));
  nor2   g0075(.a(G2104), .b(n448), .O(n449));
  nor2   g0076(.a(n449), .b(n431), .O(n450));
  inv1   g0077(.a(n450), .O(n451));
  nor2   g0078(.a(n451), .b(n447), .O(n452));
  inv1   g0079(.a(G100), .O(n453));
  nor2   g0080(.a(n429), .b(n453), .O(n454));
  inv1   g0081(.a(G136), .O(n455));
  nor2   g0082(.a(G2104), .b(n455), .O(n456));
  nor2   g0083(.a(n456), .b(G2105), .O(n457));
  inv1   g0084(.a(n457), .O(n458));
  nor2   g0085(.a(n458), .b(n454), .O(n459));
  nor2   g0086(.a(n459), .b(n452), .O(n460));
  inv1   g0087(.a(n460), .O(G162));
  inv1   g0088(.a(G114), .O(n462));
  nor2   g0089(.a(n429), .b(n462), .O(n463));
  inv1   g0090(.a(G126), .O(n464));
  nor2   g0091(.a(G2104), .b(n464), .O(n465));
  nor2   g0092(.a(n465), .b(n431), .O(n466));
  inv1   g0093(.a(n466), .O(n467));
  nor2   g0094(.a(n467), .b(n463), .O(n468));
  inv1   g0095(.a(G102), .O(n469));
  nor2   g0096(.a(n429), .b(n469), .O(n470));
  inv1   g0097(.a(G138), .O(n471));
  nor2   g0098(.a(G2104), .b(n471), .O(n472));
  nor2   g0099(.a(n472), .b(G2105), .O(n473));
  inv1   g0100(.a(n473), .O(n474));
  nor2   g0101(.a(n474), .b(n470), .O(n475));
  nor2   g0102(.a(n475), .b(n468), .O(n476));
  inv1   g0103(.a(n476), .O(G164));
  inv1   g0104(.a(G75), .O(n478));
  inv1   g0105(.a(G543), .O(n479));
  nor2   g0106(.a(n479), .b(n478), .O(n480));
  inv1   g0107(.a(G651), .O(n481));
  inv1   g0108(.a(G62), .O(n482));
  nor2   g0109(.a(G543), .b(n482), .O(n483));
  nor2   g0110(.a(n483), .b(n481), .O(n484));
  inv1   g0111(.a(n484), .O(n485));
  nor2   g0112(.a(n485), .b(n480), .O(n486));
  inv1   g0113(.a(G50), .O(n487));
  nor2   g0114(.a(n479), .b(n487), .O(n488));
  inv1   g0115(.a(G88), .O(n489));
  nor2   g0116(.a(G543), .b(n489), .O(n490));
  nor2   g0117(.a(n490), .b(G651), .O(n491));
  inv1   g0118(.a(n491), .O(n492));
  nor2   g0119(.a(n492), .b(n488), .O(n493));
  nor2   g0120(.a(n493), .b(n486), .O(G303));
  inv1   g0121(.a(G303), .O(G166));
  inv1   g0122(.a(G76), .O(n496));
  nor2   g0123(.a(n479), .b(n496), .O(n497));
  inv1   g0124(.a(G63), .O(n498));
  nor2   g0125(.a(G543), .b(n498), .O(n499));
  nor2   g0126(.a(n499), .b(n481), .O(n500));
  inv1   g0127(.a(n500), .O(n501));
  nor2   g0128(.a(n501), .b(n497), .O(n502));
  inv1   g0129(.a(G51), .O(n503));
  nor2   g0130(.a(n479), .b(n503), .O(n504));
  inv1   g0131(.a(G89), .O(n505));
  nor2   g0132(.a(G543), .b(n505), .O(n506));
  nor2   g0133(.a(n506), .b(G651), .O(n507));
  inv1   g0134(.a(n507), .O(n508));
  nor2   g0135(.a(n508), .b(n504), .O(n509));
  nor2   g0136(.a(n509), .b(n502), .O(G286));
  inv1   g0137(.a(G286), .O(G168));
  inv1   g0138(.a(G77), .O(n512));
  nor2   g0139(.a(n479), .b(n512), .O(n513));
  inv1   g0140(.a(G64), .O(n514));
  nor2   g0141(.a(G543), .b(n514), .O(n515));
  nor2   g0142(.a(n515), .b(n481), .O(n516));
  inv1   g0143(.a(n516), .O(n517));
  nor2   g0144(.a(n517), .b(n513), .O(n518));
  inv1   g0145(.a(G52), .O(n519));
  nor2   g0146(.a(n479), .b(n519), .O(n520));
  inv1   g0147(.a(G90), .O(n521));
  nor2   g0148(.a(G543), .b(n521), .O(n522));
  nor2   g0149(.a(n522), .b(G651), .O(n523));
  inv1   g0150(.a(n523), .O(n524));
  nor2   g0151(.a(n524), .b(n520), .O(n525));
  nor2   g0152(.a(n525), .b(n518), .O(G301));
  inv1   g0153(.a(G301), .O(G171));
  inv1   g0154(.a(G860), .O(n528));
  inv1   g0155(.a(G68), .O(n529));
  nor2   g0156(.a(n479), .b(n529), .O(n530));
  inv1   g0157(.a(G56), .O(n531));
  nor2   g0158(.a(G543), .b(n531), .O(n532));
  nor2   g0159(.a(n532), .b(n481), .O(n533));
  inv1   g0160(.a(n533), .O(n534));
  nor2   g0161(.a(n534), .b(n530), .O(n535));
  inv1   g0162(.a(G43), .O(n536));
  nor2   g0163(.a(n479), .b(n536), .O(n537));
  inv1   g0164(.a(G81), .O(n538));
  nor2   g0165(.a(G543), .b(n538), .O(n539));
  nor2   g0166(.a(n539), .b(G651), .O(n540));
  inv1   g0167(.a(n540), .O(n541));
  nor2   g0168(.a(n541), .b(n537), .O(n542));
  nor2   g0169(.a(n542), .b(n535), .O(n543));
  nor2   g0170(.a(n543), .b(n528), .O(n544));
  inv1   g0171(.a(n544), .O(G153));
  inv1   g0172(.a(G319), .O(n546));
  inv1   g0173(.a(G36), .O(n547));
  inv1   g0174(.a(G483), .O(n548));
  nor2   g0175(.a(n392), .b(n548), .O(n549));
  inv1   g0176(.a(n549), .O(n550));
  nor2   g0177(.a(n550), .b(n547), .O(n551));
  inv1   g0178(.a(n551), .O(n552));
  nor2   g0179(.a(n552), .b(n546), .O(n553));
  inv1   g0180(.a(n553), .O(G176));
  inv1   g0181(.a(G1), .O(n555));
  inv1   g0182(.a(G3), .O(n556));
  nor2   g0183(.a(n556), .b(n555), .O(n557));
  nor2   g0184(.a(n557), .b(n550), .O(n558));
  inv1   g0185(.a(n558), .O(n559));
  nor2   g0186(.a(n559), .b(n546), .O(n560));
  inv1   g0187(.a(n560), .O(G188));
  inv1   g0188(.a(G78), .O(n562));
  nor2   g0189(.a(n479), .b(n562), .O(n563));
  inv1   g0190(.a(G65), .O(n564));
  nor2   g0191(.a(G543), .b(n564), .O(n565));
  nor2   g0192(.a(n565), .b(n481), .O(n566));
  inv1   g0193(.a(n566), .O(n567));
  nor2   g0194(.a(n567), .b(n563), .O(n568));
  inv1   g0195(.a(G53), .O(n569));
  nor2   g0196(.a(n479), .b(n569), .O(n570));
  inv1   g0197(.a(G91), .O(n571));
  nor2   g0198(.a(G543), .b(n571), .O(n572));
  nor2   g0199(.a(n572), .b(G651), .O(n573));
  inv1   g0200(.a(n573), .O(n574));
  nor2   g0201(.a(n574), .b(n570), .O(n575));
  nor2   g0202(.a(n575), .b(n568), .O(G299));
  inv1   g0203(.a(G74), .O(n577));
  nor2   g0204(.a(n481), .b(n577), .O(n578));
  inv1   g0205(.a(G49), .O(n579));
  nor2   g0206(.a(G651), .b(n579), .O(n580));
  nor2   g0207(.a(n580), .b(n479), .O(n581));
  inv1   g0208(.a(n581), .O(n582));
  nor2   g0209(.a(n582), .b(n578), .O(n583));
  nor2   g0210(.a(G543), .b(G87), .O(n584));
  inv1   g0211(.a(n584), .O(n585));
  nor2   g0212(.a(n585), .b(G651), .O(n586));
  nor2   g0213(.a(n586), .b(n583), .O(G288));
  inv1   g0214(.a(G73), .O(n588));
  nor2   g0215(.a(n479), .b(n588), .O(n589));
  inv1   g0216(.a(G61), .O(n590));
  nor2   g0217(.a(G543), .b(n590), .O(n591));
  nor2   g0218(.a(n591), .b(n481), .O(n592));
  inv1   g0219(.a(n592), .O(n593));
  nor2   g0220(.a(n593), .b(n589), .O(n594));
  inv1   g0221(.a(G48), .O(n595));
  nor2   g0222(.a(n479), .b(n595), .O(n596));
  inv1   g0223(.a(G86), .O(n597));
  nor2   g0224(.a(G543), .b(n597), .O(n598));
  nor2   g0225(.a(n598), .b(G651), .O(n599));
  inv1   g0226(.a(n599), .O(n600));
  nor2   g0227(.a(n600), .b(n596), .O(n601));
  nor2   g0228(.a(n601), .b(n594), .O(G305));
  inv1   g0229(.a(G72), .O(n603));
  nor2   g0230(.a(n479), .b(n603), .O(n604));
  inv1   g0231(.a(G60), .O(n605));
  nor2   g0232(.a(G543), .b(n605), .O(n606));
  nor2   g0233(.a(n606), .b(n481), .O(n607));
  inv1   g0234(.a(n607), .O(n608));
  nor2   g0235(.a(n608), .b(n604), .O(n609));
  inv1   g0236(.a(G47), .O(n610));
  nor2   g0237(.a(n479), .b(n610), .O(n611));
  inv1   g0238(.a(G85), .O(n612));
  nor2   g0239(.a(G543), .b(n612), .O(n613));
  nor2   g0240(.a(n613), .b(G651), .O(n614));
  inv1   g0241(.a(n614), .O(n615));
  nor2   g0242(.a(n615), .b(n611), .O(n616));
  nor2   g0243(.a(n616), .b(n609), .O(G290));
  inv1   g0244(.a(G868), .O(n618));
  nor2   g0245(.a(G301), .b(n618), .O(n619));
  inv1   g0246(.a(G79), .O(n620));
  nor2   g0247(.a(n479), .b(n620), .O(n621));
  inv1   g0248(.a(G66), .O(n622));
  nor2   g0249(.a(G543), .b(n622), .O(n623));
  nor2   g0250(.a(n623), .b(n481), .O(n624));
  inv1   g0251(.a(n624), .O(n625));
  nor2   g0252(.a(n625), .b(n621), .O(n626));
  inv1   g0253(.a(G54), .O(n627));
  nor2   g0254(.a(n479), .b(n627), .O(n628));
  inv1   g0255(.a(G92), .O(n629));
  nor2   g0256(.a(G543), .b(n629), .O(n630));
  nor2   g0257(.a(n630), .b(G651), .O(n631));
  inv1   g0258(.a(n631), .O(n632));
  nor2   g0259(.a(n632), .b(n628), .O(n633));
  nor2   g0260(.a(n633), .b(n626), .O(n634));
  nor2   g0261(.a(n634), .b(G868), .O(n635));
  nor2   g0262(.a(n635), .b(n619), .O(G284));
  nor2   g0263(.a(G286), .b(n618), .O(n637));
  nor2   g0264(.a(G299), .b(G868), .O(n638));
  nor2   g0265(.a(n638), .b(n637), .O(G297));
  inv1   g0266(.a(G559), .O(n640));
  nor2   g0267(.a(G860), .b(n640), .O(n641));
  nor2   g0268(.a(n641), .b(n634), .O(n642));
  inv1   g0269(.a(n642), .O(G148));
  nor2   g0270(.a(n634), .b(G559), .O(n644));
  nor2   g0271(.a(n644), .b(n618), .O(n645));
  inv1   g0272(.a(n543), .O(n646));
  nor2   g0273(.a(n646), .b(G868), .O(n647));
  nor2   g0274(.a(n647), .b(n645), .O(n648));
  inv1   g0275(.a(n648), .O(G282));
  inv1   g0276(.a(G2096), .O(n650));
  inv1   g0277(.a(G111), .O(n651));
  nor2   g0278(.a(n429), .b(n651), .O(n652));
  inv1   g0279(.a(G123), .O(n653));
  nor2   g0280(.a(G2104), .b(n653), .O(n654));
  nor2   g0281(.a(n654), .b(n431), .O(n655));
  inv1   g0282(.a(n655), .O(n656));
  nor2   g0283(.a(n656), .b(n652), .O(n657));
  inv1   g0284(.a(G99), .O(n658));
  nor2   g0285(.a(n429), .b(n658), .O(n659));
  inv1   g0286(.a(G135), .O(n660));
  nor2   g0287(.a(G2104), .b(n660), .O(n661));
  nor2   g0288(.a(n661), .b(G2105), .O(n662));
  inv1   g0289(.a(n662), .O(n663));
  nor2   g0290(.a(n663), .b(n659), .O(n664));
  nor2   g0291(.a(n664), .b(n657), .O(n665));
  inv1   g0292(.a(n665), .O(n666));
  nor2   g0293(.a(n666), .b(n650), .O(n667));
  nor2   g0294(.a(n665), .b(G2096), .O(n668));
  nor2   g0295(.a(n668), .b(G2100), .O(n669));
  inv1   g0296(.a(n669), .O(n670));
  nor2   g0297(.a(n670), .b(n667), .O(n671));
  inv1   g0298(.a(n671), .O(G156));
  inv1   g0299(.a(G1341), .O(n673));
  nor2   g0300(.a(G1348), .b(n673), .O(n674));
  inv1   g0301(.a(G1348), .O(n675));
  nor2   g0302(.a(n675), .b(G1341), .O(n676));
  nor2   g0303(.a(n676), .b(n674), .O(n677));
  inv1   g0304(.a(G2427), .O(n678));
  nor2   g0305(.a(G2446), .b(G2443), .O(n679));
  inv1   g0306(.a(G2443), .O(n680));
  inv1   g0307(.a(G2446), .O(n681));
  nor2   g0308(.a(n681), .b(n680), .O(n682));
  nor2   g0309(.a(n682), .b(n679), .O(n683));
  inv1   g0310(.a(n683), .O(n684));
  nor2   g0311(.a(n684), .b(n678), .O(n685));
  nor2   g0312(.a(n683), .b(G2427), .O(n686));
  nor2   g0313(.a(n686), .b(n685), .O(n687));
  nor2   g0314(.a(G2454), .b(G2451), .O(n688));
  inv1   g0315(.a(G2451), .O(n689));
  inv1   g0316(.a(G2454), .O(n690));
  nor2   g0317(.a(n690), .b(n689), .O(n691));
  nor2   g0318(.a(n691), .b(n688), .O(n692));
  inv1   g0319(.a(n692), .O(n693));
  inv1   g0320(.a(G2430), .O(n694));
  nor2   g0321(.a(G2438), .b(G2435), .O(n695));
  inv1   g0322(.a(G2435), .O(n696));
  inv1   g0323(.a(G2438), .O(n697));
  nor2   g0324(.a(n697), .b(n696), .O(n698));
  nor2   g0325(.a(n698), .b(n695), .O(n699));
  inv1   g0326(.a(n699), .O(n700));
  nor2   g0327(.a(n700), .b(n694), .O(n701));
  nor2   g0328(.a(n699), .b(G2430), .O(n702));
  nor2   g0329(.a(n702), .b(n701), .O(n703));
  nor2   g0330(.a(n703), .b(n693), .O(n704));
  inv1   g0331(.a(n703), .O(n705));
  nor2   g0332(.a(n705), .b(n692), .O(n706));
  nor2   g0333(.a(n706), .b(n704), .O(n707));
  inv1   g0334(.a(n707), .O(n708));
  nor2   g0335(.a(n708), .b(n687), .O(n709));
  inv1   g0336(.a(n687), .O(n710));
  nor2   g0337(.a(n707), .b(n710), .O(n711));
  nor2   g0338(.a(n711), .b(n709), .O(n712));
  nor2   g0339(.a(n712), .b(n677), .O(n713));
  inv1   g0340(.a(G14), .O(n714));
  inv1   g0341(.a(n677), .O(n715));
  inv1   g0342(.a(n712), .O(n716));
  nor2   g0343(.a(n716), .b(n715), .O(n717));
  nor2   g0344(.a(n717), .b(n714), .O(n718));
  inv1   g0345(.a(n718), .O(n719));
  nor2   g0346(.a(n719), .b(n713), .O(G401));
  nor2   g0347(.a(G2100), .b(n650), .O(n721));
  inv1   g0348(.a(G2100), .O(n722));
  nor2   g0349(.a(n722), .b(G2096), .O(n723));
  nor2   g0350(.a(n723), .b(n721), .O(n724));
  inv1   g0351(.a(n724), .O(n725));
  nor2   g0352(.a(G2090), .b(G2084), .O(n726));
  nor2   g0353(.a(n726), .b(n388), .O(n727));
  inv1   g0354(.a(n727), .O(n728));
  nor2   g0355(.a(G2078), .b(G2072), .O(n729));
  nor2   g0356(.a(n729), .b(n384), .O(n730));
  inv1   g0357(.a(n730), .O(n731));
  inv1   g0358(.a(G2067), .O(n732));
  nor2   g0359(.a(G2678), .b(n732), .O(n733));
  inv1   g0360(.a(G2678), .O(n734));
  nor2   g0361(.a(n734), .b(G2067), .O(n735));
  nor2   g0362(.a(n735), .b(n733), .O(n736));
  inv1   g0363(.a(n736), .O(n737));
  nor2   g0364(.a(n737), .b(n731), .O(n738));
  nor2   g0365(.a(n736), .b(n730), .O(n739));
  nor2   g0366(.a(n739), .b(n738), .O(n740));
  nor2   g0367(.a(n740), .b(n728), .O(n741));
  inv1   g0368(.a(n740), .O(n742));
  nor2   g0369(.a(n742), .b(n727), .O(n743));
  nor2   g0370(.a(n743), .b(n741), .O(n744));
  inv1   g0371(.a(n744), .O(n745));
  nor2   g0372(.a(n745), .b(n725), .O(n746));
  nor2   g0373(.a(n744), .b(n724), .O(n747));
  nor2   g0374(.a(n747), .b(n746), .O(G227));
  nor2   g0375(.a(G1986), .b(G1981), .O(n749));
  inv1   g0376(.a(G1981), .O(n750));
  inv1   g0377(.a(G1986), .O(n751));
  nor2   g0378(.a(n751), .b(n750), .O(n752));
  nor2   g0379(.a(n752), .b(n749), .O(n753));
  inv1   g0380(.a(n753), .O(n754));
  inv1   g0381(.a(G1956), .O(n755));
  nor2   g0382(.a(G1976), .b(G1971), .O(n756));
  inv1   g0383(.a(G1971), .O(n757));
  inv1   g0384(.a(G1976), .O(n758));
  nor2   g0385(.a(n758), .b(n757), .O(n759));
  nor2   g0386(.a(n759), .b(n756), .O(n760));
  inv1   g0387(.a(n760), .O(n761));
  nor2   g0388(.a(n761), .b(n755), .O(n762));
  nor2   g0389(.a(n760), .b(G1956), .O(n763));
  nor2   g0390(.a(n763), .b(n762), .O(n764));
  nor2   g0391(.a(n764), .b(n754), .O(n765));
  inv1   g0392(.a(n764), .O(n766));
  nor2   g0393(.a(n766), .b(n753), .O(n767));
  nor2   g0394(.a(n767), .b(n765), .O(n768));
  inv1   g0395(.a(n768), .O(n769));
  inv1   g0396(.a(G2474), .O(n770));
  nor2   g0397(.a(G1966), .b(G1961), .O(n771));
  inv1   g0398(.a(G1961), .O(n772));
  inv1   g0399(.a(G1966), .O(n773));
  nor2   g0400(.a(n773), .b(n772), .O(n774));
  nor2   g0401(.a(n774), .b(n771), .O(n775));
  inv1   g0402(.a(n775), .O(n776));
  nor2   g0403(.a(n776), .b(n770), .O(n777));
  nor2   g0404(.a(n775), .b(G2474), .O(n778));
  nor2   g0405(.a(n778), .b(n777), .O(n779));
  inv1   g0406(.a(n779), .O(n780));
  inv1   g0407(.a(G1991), .O(n781));
  nor2   g0408(.a(G1996), .b(n781), .O(n782));
  inv1   g0409(.a(G1996), .O(n783));
  nor2   g0410(.a(n783), .b(G1991), .O(n784));
  nor2   g0411(.a(n784), .b(n782), .O(n785));
  nor2   g0412(.a(n785), .b(n780), .O(n786));
  inv1   g0413(.a(n785), .O(n787));
  nor2   g0414(.a(n787), .b(n779), .O(n788));
  nor2   g0415(.a(n788), .b(n786), .O(n789));
  inv1   g0416(.a(n789), .O(n790));
  nor2   g0417(.a(n790), .b(n769), .O(n791));
  nor2   g0418(.a(n789), .b(n768), .O(n792));
  nor2   g0419(.a(n792), .b(n791), .O(G229));
  nor2   g0420(.a(G29), .b(G26), .O(n794));
  inv1   g0421(.a(G29), .O(n795));
  inv1   g0422(.a(G116), .O(n796));
  nor2   g0423(.a(n429), .b(n796), .O(n797));
  inv1   g0424(.a(G128), .O(n798));
  nor2   g0425(.a(G2104), .b(n798), .O(n799));
  nor2   g0426(.a(n799), .b(n431), .O(n800));
  inv1   g0427(.a(n800), .O(n801));
  nor2   g0428(.a(n801), .b(n797), .O(n802));
  inv1   g0429(.a(G104), .O(n803));
  nor2   g0430(.a(n429), .b(n803), .O(n804));
  inv1   g0431(.a(G140), .O(n805));
  nor2   g0432(.a(G2104), .b(n805), .O(n806));
  nor2   g0433(.a(n806), .b(G2105), .O(n807));
  inv1   g0434(.a(n807), .O(n808));
  nor2   g0435(.a(n808), .b(n804), .O(n809));
  nor2   g0436(.a(n809), .b(n802), .O(n810));
  nor2   g0437(.a(n810), .b(n795), .O(n811));
  nor2   g0438(.a(n811), .b(n794), .O(n812));
  inv1   g0439(.a(n812), .O(n813));
  nor2   g0440(.a(n813), .b(n732), .O(n814));
  nor2   g0441(.a(G35), .b(G29), .O(n815));
  nor2   g0442(.a(n460), .b(n795), .O(n816));
  nor2   g0443(.a(n816), .b(n815), .O(n817));
  nor2   g0444(.a(n817), .b(G2090), .O(n818));
  nor2   g0445(.a(G16), .b(G6), .O(n819));
  inv1   g0446(.a(G16), .O(n820));
  nor2   g0447(.a(G305), .b(n820), .O(n821));
  nor2   g0448(.a(n821), .b(n819), .O(n822));
  inv1   g0449(.a(n822), .O(n823));
  nor2   g0450(.a(n823), .b(n750), .O(n824));
  nor2   g0451(.a(n824), .b(n818), .O(n825));
  inv1   g0452(.a(n825), .O(n826));
  nor2   g0453(.a(n826), .b(n814), .O(n827));
  inv1   g0454(.a(n827), .O(n828));
  inv1   g0455(.a(n817), .O(n829));
  nor2   g0456(.a(n829), .b(n387), .O(n830));
  nor2   g0457(.a(G16), .b(G4), .O(n831));
  nor2   g0458(.a(n634), .b(n820), .O(n832));
  nor2   g0459(.a(n832), .b(n831), .O(n833));
  inv1   g0460(.a(n833), .O(n834));
  nor2   g0461(.a(n834), .b(n675), .O(n835));
  nor2   g0462(.a(n835), .b(n830), .O(n836));
  inv1   g0463(.a(n836), .O(n837));
  nor2   g0464(.a(G19), .b(G16), .O(n838));
  nor2   g0465(.a(n543), .b(n820), .O(n839));
  nor2   g0466(.a(n839), .b(n838), .O(n840));
  nor2   g0467(.a(n840), .b(G1341), .O(n841));
  nor2   g0468(.a(G34), .b(G29), .O(n842));
  nor2   g0469(.a(n444), .b(n795), .O(n843));
  nor2   g0470(.a(n843), .b(n842), .O(n844));
  inv1   g0471(.a(n844), .O(n845));
  nor2   g0472(.a(n845), .b(n386), .O(n846));
  nor2   g0473(.a(n846), .b(n841), .O(n847));
  inv1   g0474(.a(n847), .O(n848));
  nor2   g0475(.a(n848), .b(n837), .O(n849));
  inv1   g0476(.a(n849), .O(n850));
  nor2   g0477(.a(G33), .b(G29), .O(n851));
  inv1   g0478(.a(G115), .O(n852));
  nor2   g0479(.a(n429), .b(n852), .O(n853));
  inv1   g0480(.a(G127), .O(n854));
  nor2   g0481(.a(G2104), .b(n854), .O(n855));
  nor2   g0482(.a(n855), .b(n431), .O(n856));
  inv1   g0483(.a(n856), .O(n857));
  nor2   g0484(.a(n857), .b(n853), .O(n858));
  inv1   g0485(.a(G103), .O(n859));
  nor2   g0486(.a(n429), .b(n859), .O(n860));
  inv1   g0487(.a(G139), .O(n861));
  nor2   g0488(.a(G2104), .b(n861), .O(n862));
  nor2   g0489(.a(n862), .b(G2105), .O(n863));
  inv1   g0490(.a(n863), .O(n864));
  nor2   g0491(.a(n864), .b(n860), .O(n865));
  nor2   g0492(.a(n865), .b(n858), .O(n866));
  nor2   g0493(.a(n866), .b(n795), .O(n867));
  nor2   g0494(.a(n867), .b(n851), .O(n868));
  inv1   g0495(.a(n868), .O(n869));
  nor2   g0496(.a(n869), .b(n382), .O(n870));
  nor2   g0497(.a(n812), .b(G2067), .O(n871));
  nor2   g0498(.a(n871), .b(n870), .O(n872));
  inv1   g0499(.a(n872), .O(n873));
  nor2   g0500(.a(n822), .b(G1981), .O(n874));
  inv1   g0501(.a(n840), .O(n875));
  nor2   g0502(.a(n875), .b(n673), .O(n876));
  nor2   g0503(.a(n876), .b(n874), .O(n877));
  inv1   g0504(.a(n877), .O(n878));
  nor2   g0505(.a(n878), .b(n873), .O(n879));
  inv1   g0506(.a(n879), .O(n880));
  nor2   g0507(.a(n880), .b(n850), .O(n881));
  inv1   g0508(.a(n881), .O(n882));
  nor2   g0509(.a(n882), .b(n828), .O(n883));
  inv1   g0510(.a(n883), .O(n884));
  nor2   g0511(.a(G23), .b(G16), .O(n885));
  nor2   g0512(.a(G288), .b(n820), .O(n886));
  nor2   g0513(.a(n886), .b(n885), .O(n887));
  nor2   g0514(.a(n887), .b(n758), .O(n888));
  inv1   g0515(.a(n887), .O(n889));
  nor2   g0516(.a(n889), .b(G1976), .O(n890));
  nor2   g0517(.a(n890), .b(n888), .O(n891));
  nor2   g0518(.a(G29), .b(G27), .O(n892));
  nor2   g0519(.a(n476), .b(n795), .O(n893));
  nor2   g0520(.a(n893), .b(n892), .O(n894));
  nor2   g0521(.a(n894), .b(n383), .O(n895));
  inv1   g0522(.a(n894), .O(n896));
  nor2   g0523(.a(n896), .b(G2078), .O(n897));
  nor2   g0524(.a(n897), .b(n895), .O(n898));
  nor2   g0525(.a(G29), .b(G25), .O(n899));
  inv1   g0526(.a(G107), .O(n900));
  nor2   g0527(.a(n429), .b(n900), .O(n901));
  inv1   g0528(.a(G119), .O(n902));
  nor2   g0529(.a(G2104), .b(n902), .O(n903));
  nor2   g0530(.a(n903), .b(n431), .O(n904));
  inv1   g0531(.a(n904), .O(n905));
  nor2   g0532(.a(n905), .b(n901), .O(n906));
  inv1   g0533(.a(G95), .O(n907));
  nor2   g0534(.a(n429), .b(n907), .O(n908));
  inv1   g0535(.a(G131), .O(n909));
  nor2   g0536(.a(G2104), .b(n909), .O(n910));
  nor2   g0537(.a(n910), .b(G2105), .O(n911));
  inv1   g0538(.a(n911), .O(n912));
  nor2   g0539(.a(n912), .b(n908), .O(n913));
  nor2   g0540(.a(n913), .b(n906), .O(n914));
  nor2   g0541(.a(n914), .b(n795), .O(n915));
  nor2   g0542(.a(n915), .b(n899), .O(n916));
  nor2   g0543(.a(n916), .b(n781), .O(n917));
  inv1   g0544(.a(n916), .O(n918));
  nor2   g0545(.a(n918), .b(G1991), .O(n919));
  nor2   g0546(.a(n919), .b(n917), .O(n920));
  nor2   g0547(.a(n920), .b(n898), .O(n921));
  inv1   g0548(.a(n921), .O(n922));
  nor2   g0549(.a(n922), .b(n891), .O(n923));
  inv1   g0550(.a(n923), .O(n924));
  nor2   g0551(.a(n868), .b(G2072), .O(n925));
  nor2   g0552(.a(n665), .b(n795), .O(n926));
  inv1   g0553(.a(G11), .O(n927));
  nor2   g0554(.a(G29), .b(G28), .O(n928));
  nor2   g0555(.a(n928), .b(n927), .O(n929));
  inv1   g0556(.a(n929), .O(n930));
  nor2   g0557(.a(n930), .b(n926), .O(n931));
  inv1   g0558(.a(n931), .O(n932));
  nor2   g0559(.a(n932), .b(n925), .O(n933));
  inv1   g0560(.a(n933), .O(n934));
  nor2   g0561(.a(G32), .b(G29), .O(n935));
  inv1   g0562(.a(G117), .O(n936));
  nor2   g0563(.a(n429), .b(n936), .O(n937));
  inv1   g0564(.a(G129), .O(n938));
  nor2   g0565(.a(G2104), .b(n938), .O(n939));
  nor2   g0566(.a(n939), .b(n431), .O(n940));
  inv1   g0567(.a(n940), .O(n941));
  nor2   g0568(.a(n941), .b(n937), .O(n942));
  inv1   g0569(.a(G105), .O(n943));
  nor2   g0570(.a(n429), .b(n943), .O(n944));
  inv1   g0571(.a(G141), .O(n945));
  nor2   g0572(.a(G2104), .b(n945), .O(n946));
  nor2   g0573(.a(n946), .b(G2105), .O(n947));
  inv1   g0574(.a(n947), .O(n948));
  nor2   g0575(.a(n948), .b(n944), .O(n949));
  nor2   g0576(.a(n949), .b(n942), .O(n950));
  nor2   g0577(.a(n950), .b(n795), .O(n951));
  nor2   g0578(.a(n951), .b(n935), .O(n952));
  inv1   g0579(.a(n952), .O(n953));
  nor2   g0580(.a(n953), .b(n783), .O(n954));
  nor2   g0581(.a(n833), .b(G1348), .O(n955));
  nor2   g0582(.a(n955), .b(n954), .O(n956));
  inv1   g0583(.a(n956), .O(n957));
  nor2   g0584(.a(n957), .b(n934), .O(n958));
  inv1   g0585(.a(n958), .O(n959));
  nor2   g0586(.a(G22), .b(G16), .O(n960));
  nor2   g0587(.a(G303), .b(n820), .O(n961));
  nor2   g0588(.a(n961), .b(n960), .O(n962));
  nor2   g0589(.a(n962), .b(n757), .O(n963));
  inv1   g0590(.a(n962), .O(n964));
  nor2   g0591(.a(n964), .b(G1971), .O(n965));
  nor2   g0592(.a(n965), .b(n963), .O(n966));
  nor2   g0593(.a(G16), .b(G5), .O(n967));
  nor2   g0594(.a(G301), .b(n820), .O(n968));
  nor2   g0595(.a(n968), .b(n967), .O(n969));
  nor2   g0596(.a(n969), .b(n772), .O(n970));
  inv1   g0597(.a(n969), .O(n971));
  nor2   g0598(.a(n971), .b(G1961), .O(n972));
  nor2   g0599(.a(n972), .b(n970), .O(n973));
  nor2   g0600(.a(n973), .b(n966), .O(n974));
  inv1   g0601(.a(n974), .O(n975));
  nor2   g0602(.a(n975), .b(n959), .O(n976));
  inv1   g0603(.a(n976), .O(n977));
  nor2   g0604(.a(G24), .b(G16), .O(n978));
  nor2   g0605(.a(G290), .b(n820), .O(n979));
  nor2   g0606(.a(n979), .b(n978), .O(n980));
  inv1   g0607(.a(n980), .O(n981));
  nor2   g0608(.a(n981), .b(n751), .O(n982));
  nor2   g0609(.a(n952), .b(G1996), .O(n983));
  nor2   g0610(.a(n983), .b(n982), .O(n984));
  inv1   g0611(.a(n984), .O(n985));
  nor2   g0612(.a(n844), .b(G2084), .O(n986));
  nor2   g0613(.a(G21), .b(G16), .O(n987));
  nor2   g0614(.a(G286), .b(n820), .O(n988));
  nor2   g0615(.a(n988), .b(n987), .O(n989));
  inv1   g0616(.a(n989), .O(n990));
  nor2   g0617(.a(n990), .b(n773), .O(n991));
  nor2   g0618(.a(n991), .b(n986), .O(n992));
  inv1   g0619(.a(n992), .O(n993));
  nor2   g0620(.a(n993), .b(n985), .O(n994));
  inv1   g0621(.a(n994), .O(n995));
  nor2   g0622(.a(n980), .b(G1986), .O(n996));
  nor2   g0623(.a(G20), .b(G16), .O(n997));
  nor2   g0624(.a(G299), .b(n820), .O(n998));
  nor2   g0625(.a(n998), .b(n997), .O(n999));
  inv1   g0626(.a(n999), .O(n1000));
  nor2   g0627(.a(n1000), .b(n755), .O(n1001));
  nor2   g0628(.a(n1001), .b(n996), .O(n1002));
  inv1   g0629(.a(n1002), .O(n1003));
  nor2   g0630(.a(n989), .b(G1966), .O(n1004));
  nor2   g0631(.a(n999), .b(G1956), .O(n1005));
  nor2   g0632(.a(n1005), .b(n1004), .O(n1006));
  inv1   g0633(.a(n1006), .O(n1007));
  nor2   g0634(.a(n1007), .b(n1003), .O(n1008));
  inv1   g0635(.a(n1008), .O(n1009));
  nor2   g0636(.a(n1009), .b(n995), .O(n1010));
  inv1   g0637(.a(n1010), .O(n1011));
  nor2   g0638(.a(n1011), .b(n977), .O(n1012));
  inv1   g0639(.a(n1012), .O(n1013));
  nor2   g0640(.a(n1013), .b(n924), .O(n1014));
  inv1   g0641(.a(n1014), .O(n1015));
  nor2   g0642(.a(n1015), .b(n884), .O(G311));
  inv1   g0643(.a(G311), .O(G150));
  inv1   g0644(.a(n641), .O(n1018));
  nor2   g0645(.a(n1018), .b(n634), .O(n1019));
  nor2   g0646(.a(n1019), .b(n544), .O(n1020));
  inv1   g0647(.a(G80), .O(n1021));
  nor2   g0648(.a(n479), .b(n1021), .O(n1022));
  inv1   g0649(.a(G67), .O(n1023));
  nor2   g0650(.a(G543), .b(n1023), .O(n1024));
  nor2   g0651(.a(n1024), .b(n481), .O(n1025));
  inv1   g0652(.a(n1025), .O(n1026));
  nor2   g0653(.a(n1026), .b(n1022), .O(n1027));
  inv1   g0654(.a(G55), .O(n1028));
  nor2   g0655(.a(n479), .b(n1028), .O(n1029));
  inv1   g0656(.a(G93), .O(n1030));
  nor2   g0657(.a(G543), .b(n1030), .O(n1031));
  nor2   g0658(.a(n1031), .b(G651), .O(n1032));
  inv1   g0659(.a(n1032), .O(n1033));
  nor2   g0660(.a(n1033), .b(n1029), .O(n1034));
  nor2   g0661(.a(n1034), .b(n1027), .O(n1035));
  nor2   g0662(.a(n1035), .b(n543), .O(n1036));
  inv1   g0663(.a(n1035), .O(n1037));
  nor2   g0664(.a(n1037), .b(n646), .O(n1038));
  nor2   g0665(.a(n1038), .b(n1036), .O(n1039));
  nor2   g0666(.a(n1039), .b(n1020), .O(n1040));
  inv1   g0667(.a(n1020), .O(n1041));
  inv1   g0668(.a(n1039), .O(n1042));
  nor2   g0669(.a(n1042), .b(n1041), .O(n1043));
  nor2   g0670(.a(n1043), .b(n1040), .O(G145));
  nor2   g0671(.a(n460), .b(G160), .O(n1045));
  nor2   g0672(.a(G162), .b(n444), .O(n1046));
  nor2   g0673(.a(n1046), .b(n1045), .O(n1047));
  inv1   g0674(.a(n1047), .O(n1048));
  nor2   g0675(.a(n1048), .b(n666), .O(n1049));
  nor2   g0676(.a(n1047), .b(n665), .O(n1050));
  nor2   g0677(.a(n1050), .b(n1049), .O(n1051));
  inv1   g0678(.a(n1051), .O(n1052));
  inv1   g0679(.a(n950), .O(n1053));
  nor2   g0680(.a(n1053), .b(n810), .O(n1054));
  inv1   g0681(.a(n810), .O(n1055));
  nor2   g0682(.a(n950), .b(n1055), .O(n1056));
  nor2   g0683(.a(n1056), .b(n1054), .O(n1057));
  inv1   g0684(.a(n1057), .O(n1058));
  inv1   g0685(.a(G118), .O(n1059));
  nor2   g0686(.a(n429), .b(n1059), .O(n1060));
  inv1   g0687(.a(G130), .O(n1061));
  nor2   g0688(.a(G2104), .b(n1061), .O(n1062));
  nor2   g0689(.a(n1062), .b(n431), .O(n1063));
  inv1   g0690(.a(n1063), .O(n1064));
  nor2   g0691(.a(n1064), .b(n1060), .O(n1065));
  inv1   g0692(.a(G106), .O(n1066));
  nor2   g0693(.a(n429), .b(n1066), .O(n1067));
  inv1   g0694(.a(G142), .O(n1068));
  nor2   g0695(.a(G2104), .b(n1068), .O(n1069));
  nor2   g0696(.a(n1069), .b(G2105), .O(n1070));
  inv1   g0697(.a(n1070), .O(n1071));
  nor2   g0698(.a(n1071), .b(n1067), .O(n1072));
  nor2   g0699(.a(n1072), .b(n1065), .O(n1073));
  inv1   g0700(.a(n1073), .O(n1074));
  inv1   g0701(.a(n866), .O(n1075));
  nor2   g0702(.a(n914), .b(G164), .O(n1076));
  inv1   g0703(.a(n914), .O(n1077));
  nor2   g0704(.a(n1077), .b(n476), .O(n1078));
  nor2   g0705(.a(n1078), .b(n1076), .O(n1079));
  inv1   g0706(.a(n1079), .O(n1080));
  nor2   g0707(.a(n1080), .b(n1075), .O(n1081));
  nor2   g0708(.a(n1079), .b(n866), .O(n1082));
  nor2   g0709(.a(n1082), .b(n1081), .O(n1083));
  nor2   g0710(.a(n1083), .b(n1074), .O(n1084));
  inv1   g0711(.a(n1083), .O(n1085));
  nor2   g0712(.a(n1085), .b(n1073), .O(n1086));
  nor2   g0713(.a(n1086), .b(n1084), .O(n1087));
  inv1   g0714(.a(n1087), .O(n1088));
  nor2   g0715(.a(n1088), .b(n1058), .O(n1089));
  nor2   g0716(.a(n1087), .b(n1057), .O(n1090));
  nor2   g0717(.a(n1090), .b(n1089), .O(n1091));
  inv1   g0718(.a(n1091), .O(n1092));
  nor2   g0719(.a(n1092), .b(n1052), .O(n1093));
  nor2   g0720(.a(n1091), .b(n1051), .O(n1094));
  nor2   g0721(.a(n1094), .b(G37), .O(n1095));
  inv1   g0722(.a(n1095), .O(n1096));
  nor2   g0723(.a(n1096), .b(n1093), .O(G395));
  nor2   g0724(.a(G305), .b(G166), .O(n1098));
  inv1   g0725(.a(G305), .O(n1099));
  nor2   g0726(.a(n1099), .b(G303), .O(n1100));
  nor2   g0727(.a(n1100), .b(n1098), .O(n1101));
  inv1   g0728(.a(n1101), .O(n1102));
  inv1   g0729(.a(G290), .O(n1103));
  nor2   g0730(.a(n1103), .b(G288), .O(n1104));
  inv1   g0731(.a(G288), .O(n1105));
  nor2   g0732(.a(G290), .b(n1105), .O(n1106));
  nor2   g0733(.a(n1106), .b(n1104), .O(n1107));
  inv1   g0734(.a(n1107), .O(n1108));
  nor2   g0735(.a(n1108), .b(n1102), .O(n1109));
  nor2   g0736(.a(n1107), .b(n1101), .O(n1110));
  nor2   g0737(.a(n1110), .b(n1109), .O(n1111));
  inv1   g0738(.a(n1111), .O(n1112));
  inv1   g0739(.a(n644), .O(n1113));
  nor2   g0740(.a(n1039), .b(G299), .O(n1114));
  inv1   g0741(.a(G299), .O(n1115));
  nor2   g0742(.a(n1042), .b(n1115), .O(n1116));
  nor2   g0743(.a(n1116), .b(n1114), .O(n1117));
  nor2   g0744(.a(n1117), .b(n1113), .O(n1118));
  inv1   g0745(.a(n634), .O(n1119));
  nor2   g0746(.a(n1117), .b(n1119), .O(n1120));
  inv1   g0747(.a(n1117), .O(n1121));
  nor2   g0748(.a(n1121), .b(n634), .O(n1122));
  nor2   g0749(.a(n1122), .b(n1120), .O(n1123));
  nor2   g0750(.a(n1123), .b(n644), .O(n1124));
  nor2   g0751(.a(n1124), .b(n1118), .O(n1125));
  nor2   g0752(.a(n1125), .b(n1112), .O(n1126));
  inv1   g0753(.a(n1125), .O(n1127));
  nor2   g0754(.a(n1127), .b(n1111), .O(n1128));
  nor2   g0755(.a(n1128), .b(n1126), .O(n1129));
  nor2   g0756(.a(n1129), .b(n618), .O(n1130));
  nor2   g0757(.a(n1037), .b(G868), .O(n1131));
  nor2   g0758(.a(n1131), .b(n1130), .O(n1132));
  inv1   g0759(.a(n1132), .O(G295));
  inv1   g0760(.a(n1123), .O(n1134));
  nor2   g0761(.a(G301), .b(G168), .O(n1135));
  nor2   g0762(.a(G171), .b(G286), .O(n1136));
  nor2   g0763(.a(n1136), .b(n1135), .O(n1137));
  inv1   g0764(.a(n1137), .O(n1138));
  nor2   g0765(.a(n1138), .b(n1134), .O(n1139));
  nor2   g0766(.a(n1137), .b(n1123), .O(n1140));
  nor2   g0767(.a(n1140), .b(n1139), .O(n1141));
  nor2   g0768(.a(n1141), .b(n1112), .O(n1142));
  inv1   g0769(.a(n1141), .O(n1143));
  nor2   g0770(.a(n1143), .b(n1111), .O(n1144));
  nor2   g0771(.a(n1144), .b(G37), .O(n1145));
  inv1   g0772(.a(n1145), .O(n1146));
  nor2   g0773(.a(n1146), .b(n1142), .O(G397));
  nor2   g0774(.a(G164), .b(G1384), .O(n1148));
  inv1   g0775(.a(n1148), .O(n1149));
  inv1   g0776(.a(G40), .O(n1150));
  nor2   g0777(.a(n444), .b(n1150), .O(n1151));
  inv1   g0778(.a(n1151), .O(n1152));
  nor2   g0779(.a(n1152), .b(n1149), .O(n1153));
  nor2   g0780(.a(n1153), .b(n773), .O(n1154));
  inv1   g0781(.a(G8), .O(n1155));
  inv1   g0782(.a(n1153), .O(n1156));
  nor2   g0783(.a(n1156), .b(n386), .O(n1157));
  nor2   g0784(.a(n1157), .b(n1155), .O(n1158));
  inv1   g0785(.a(n1158), .O(n1159));
  nor2   g0786(.a(n1159), .b(n1154), .O(n1160));
  inv1   g0787(.a(n1160), .O(n1161));
  nor2   g0788(.a(n1161), .b(G286), .O(n1162));
  nor2   g0789(.a(G168), .b(n1155), .O(n1163));
  inv1   g0790(.a(n1163), .O(n1164));
  nor2   g0791(.a(n1164), .b(n1160), .O(n1165));
  nor2   g0792(.a(n1165), .b(n1162), .O(n1166));
  inv1   g0793(.a(n1166), .O(n1167));
  nor2   g0794(.a(n1153), .b(n757), .O(n1168));
  nor2   g0795(.a(n1156), .b(n387), .O(n1169));
  nor2   g0796(.a(n1169), .b(n1155), .O(n1170));
  inv1   g0797(.a(n1170), .O(n1171));
  nor2   g0798(.a(n1171), .b(n1168), .O(n1172));
  nor2   g0799(.a(G166), .b(n1155), .O(n1173));
  inv1   g0800(.a(n1173), .O(n1174));
  nor2   g0801(.a(n1174), .b(n1172), .O(n1175));
  inv1   g0802(.a(n1172), .O(n1176));
  nor2   g0803(.a(n1176), .b(G303), .O(n1177));
  nor2   g0804(.a(n1177), .b(n1175), .O(n1178));
  inv1   g0805(.a(n1178), .O(n1179));
  nor2   g0806(.a(n1153), .b(n772), .O(n1180));
  nor2   g0807(.a(n1156), .b(n383), .O(n1181));
  nor2   g0808(.a(n1181), .b(n1180), .O(n1182));
  inv1   g0809(.a(n1182), .O(n1183));
  nor2   g0810(.a(n1183), .b(G301), .O(n1184));
  inv1   g0811(.a(n1184), .O(n1185));
  nor2   g0812(.a(G1981), .b(n1155), .O(n1186));
  inv1   g0813(.a(n1186), .O(n1187));
  nor2   g0814(.a(n1187), .b(G305), .O(n1188));
  inv1   g0815(.a(n1188), .O(n1189));
  nor2   g0816(.a(n1189), .b(n1153), .O(n1190));
  nor2   g0817(.a(n758), .b(n1155), .O(n1191));
  inv1   g0818(.a(n1191), .O(n1192));
  nor2   g0819(.a(n1192), .b(n1105), .O(n1193));
  inv1   g0820(.a(n1193), .O(n1194));
  nor2   g0821(.a(n1194), .b(n1153), .O(n1195));
  nor2   g0822(.a(n1195), .b(n1190), .O(n1196));
  inv1   g0823(.a(n1196), .O(n1197));
  nor2   g0824(.a(n750), .b(n1155), .O(n1198));
  inv1   g0825(.a(n1198), .O(n1199));
  nor2   g0826(.a(n1199), .b(n1099), .O(n1200));
  inv1   g0827(.a(n1200), .O(n1201));
  nor2   g0828(.a(n1201), .b(n1153), .O(n1202));
  nor2   g0829(.a(G1976), .b(n1155), .O(n1203));
  inv1   g0830(.a(n1203), .O(n1204));
  nor2   g0831(.a(n1204), .b(G288), .O(n1205));
  inv1   g0832(.a(n1205), .O(n1206));
  nor2   g0833(.a(n1206), .b(n1153), .O(n1207));
  nor2   g0834(.a(n1207), .b(n1202), .O(n1208));
  inv1   g0835(.a(n1208), .O(n1209));
  nor2   g0836(.a(n1209), .b(n1197), .O(n1210));
  inv1   g0837(.a(n1210), .O(n1211));
  nor2   g0838(.a(n1211), .b(n1185), .O(n1212));
  inv1   g0839(.a(n1212), .O(n1213));
  nor2   g0840(.a(n1213), .b(n1179), .O(n1214));
  inv1   g0841(.a(n1214), .O(n1215));
  nor2   g0842(.a(n1215), .b(n1167), .O(n1216));
  nor2   g0843(.a(n1182), .b(G171), .O(n1217));
  nor2   g0844(.a(n1217), .b(n1184), .O(n1218));
  inv1   g0845(.a(n1218), .O(n1219));
  nor2   g0846(.a(n1153), .b(n755), .O(n1220));
  nor2   g0847(.a(n1156), .b(n382), .O(n1221));
  nor2   g0848(.a(n1221), .b(n1220), .O(n1222));
  nor2   g0849(.a(n1222), .b(n1115), .O(n1223));
  nor2   g0850(.a(n1223), .b(n1211), .O(n1224));
  inv1   g0851(.a(n1224), .O(n1225));
  nor2   g0852(.a(n1225), .b(n1219), .O(n1226));
  inv1   g0853(.a(n1226), .O(n1227));
  nor2   g0854(.a(n1227), .b(n1179), .O(n1228));
  inv1   g0855(.a(n1228), .O(n1229));
  nor2   g0856(.a(n1153), .b(n675), .O(n1230));
  nor2   g0857(.a(n1156), .b(n732), .O(n1231));
  nor2   g0858(.a(n1231), .b(n1230), .O(n1232));
  nor2   g0859(.a(n1232), .b(n1119), .O(n1233));
  nor2   g0860(.a(n1153), .b(n673), .O(n1234));
  nor2   g0861(.a(n1156), .b(n783), .O(n1235));
  nor2   g0862(.a(n1235), .b(n543), .O(n1236));
  inv1   g0863(.a(n1236), .O(n1237));
  nor2   g0864(.a(n1237), .b(n1234), .O(n1238));
  inv1   g0865(.a(n1238), .O(n1239));
  nor2   g0866(.a(n1239), .b(n1233), .O(n1240));
  inv1   g0867(.a(n1222), .O(n1241));
  nor2   g0868(.a(n1241), .b(G299), .O(n1242));
  inv1   g0869(.a(n1232), .O(n1243));
  nor2   g0870(.a(n1243), .b(n634), .O(n1244));
  nor2   g0871(.a(n1244), .b(n1242), .O(n1245));
  inv1   g0872(.a(n1245), .O(n1246));
  nor2   g0873(.a(n1246), .b(n1240), .O(n1247));
  nor2   g0874(.a(n1247), .b(n1167), .O(n1248));
  inv1   g0875(.a(n1248), .O(n1249));
  nor2   g0876(.a(n1249), .b(n1229), .O(n1250));
  inv1   g0877(.a(n1162), .O(n1251));
  nor2   g0878(.a(n1211), .b(n1251), .O(n1252));
  inv1   g0879(.a(n1252), .O(n1253));
  nor2   g0880(.a(n1253), .b(n1179), .O(n1254));
  inv1   g0881(.a(n1177), .O(n1255));
  nor2   g0882(.a(n1211), .b(n1255), .O(n1256));
  inv1   g0883(.a(n1207), .O(n1257));
  nor2   g0884(.a(n1257), .b(n1202), .O(n1258));
  nor2   g0885(.a(n1258), .b(n1190), .O(n1259));
  inv1   g0886(.a(n1259), .O(n1260));
  nor2   g0887(.a(n1260), .b(n1256), .O(n1261));
  inv1   g0888(.a(n1261), .O(n1262));
  nor2   g0889(.a(n1262), .b(n1254), .O(n1263));
  inv1   g0890(.a(n1263), .O(n1264));
  nor2   g0891(.a(n1264), .b(n1250), .O(n1265));
  inv1   g0892(.a(n1265), .O(n1266));
  nor2   g0893(.a(n1266), .b(n1216), .O(n1267));
  nor2   g0894(.a(n1152), .b(n1148), .O(n1268));
  inv1   g0895(.a(n1268), .O(n1269));
  nor2   g0896(.a(n1055), .b(n732), .O(n1270));
  inv1   g0897(.a(n1270), .O(n1271));
  nor2   g0898(.a(n1271), .b(n1269), .O(n1272));
  nor2   g0899(.a(n950), .b(G1996), .O(n1273));
  inv1   g0900(.a(n1273), .O(n1274));
  nor2   g0901(.a(n1274), .b(n1269), .O(n1275));
  nor2   g0902(.a(n1275), .b(n1272), .O(n1276));
  inv1   g0903(.a(n1276), .O(n1277));
  nor2   g0904(.a(n1103), .b(n751), .O(n1278));
  inv1   g0905(.a(n1278), .O(n1279));
  nor2   g0906(.a(n1279), .b(n1269), .O(n1280));
  nor2   g0907(.a(n1077), .b(n781), .O(n1281));
  inv1   g0908(.a(n1281), .O(n1282));
  nor2   g0909(.a(n1282), .b(n1269), .O(n1283));
  nor2   g0910(.a(n1283), .b(n1280), .O(n1284));
  inv1   g0911(.a(n1284), .O(n1285));
  nor2   g0912(.a(n1285), .b(n1277), .O(n1286));
  inv1   g0913(.a(n1286), .O(n1287));
  nor2   g0914(.a(G290), .b(G1986), .O(n1288));
  inv1   g0915(.a(n1288), .O(n1289));
  nor2   g0916(.a(n1289), .b(n1269), .O(n1290));
  nor2   g0917(.a(n914), .b(G1991), .O(n1291));
  inv1   g0918(.a(n1291), .O(n1292));
  nor2   g0919(.a(n1292), .b(n1269), .O(n1293));
  nor2   g0920(.a(n1293), .b(n1290), .O(n1294));
  inv1   g0921(.a(n1294), .O(n1295));
  nor2   g0922(.a(n810), .b(G2067), .O(n1296));
  inv1   g0923(.a(n1296), .O(n1297));
  nor2   g0924(.a(n1297), .b(n1269), .O(n1298));
  nor2   g0925(.a(n1053), .b(n783), .O(n1299));
  inv1   g0926(.a(n1299), .O(n1300));
  nor2   g0927(.a(n1300), .b(n1269), .O(n1301));
  nor2   g0928(.a(n1301), .b(n1298), .O(n1302));
  inv1   g0929(.a(n1302), .O(n1303));
  nor2   g0930(.a(n1303), .b(n1295), .O(n1304));
  inv1   g0931(.a(n1304), .O(n1305));
  nor2   g0932(.a(n1305), .b(n1287), .O(n1306));
  inv1   g0933(.a(n1306), .O(n1307));
  nor2   g0934(.a(n1307), .b(n1267), .O(n1308));
  nor2   g0935(.a(n1077), .b(n781), .O(n1309));
  nor2   g0936(.a(n1301), .b(n1294), .O(n1310));
  inv1   g0937(.a(n1310), .O(n1311));
  nor2   g0938(.a(n1311), .b(n1309), .O(n1312));
  nor2   g0939(.a(n1312), .b(n1275), .O(n1313));
  nor2   g0940(.a(n1313), .b(n1272), .O(n1314));
  nor2   g0941(.a(n1314), .b(n1298), .O(n1315));
  inv1   g0942(.a(n1315), .O(n1316));
  nor2   g0943(.a(n1316), .b(n1308), .O(n1317));
  inv1   g0944(.a(n1317), .O(G329));
  nor2   g0945(.a(G227), .b(n546), .O(n1320));
  inv1   g0946(.a(n1320), .O(n1321));
  nor2   g0947(.a(n1321), .b(G229), .O(n1322));
  inv1   g0948(.a(n1322), .O(n1323));
  nor2   g0949(.a(n1323), .b(G401), .O(n1324));
  inv1   g0950(.a(n1324), .O(n1325));
  nor2   g0951(.a(n1325), .b(G395), .O(n1326));
  inv1   g0952(.a(n1326), .O(n1327));
  nor2   g0953(.a(n1327), .b(G397), .O(G308));
  inv1   g0954(.a(G308), .O(G225));
  zero   g0955(.O(G231));
  buffer g0956(.a(ING169 ), .O(G169));
  buffer g0957(.a(ING174 ), .O(G174));
  buffer g0958(.a(ING177 ), .O(G177));
  buffer g0959(.a(ING178 ), .O(G178));
  buffer g0960(.a(ING179 ), .O(G179));
  buffer g0961(.a(ING180 ), .O(G180));
  buffer g0962(.a(ING181 ), .O(G181));
  buffer g0963(.a(ING182 ), .O(G182));
  buffer g0964(.a(ING183 ), .O(G183));
  buffer g0965(.a(ING184 ), .O(G184));
  buffer g0966(.a(ING185 ), .O(G185));
  buffer g0967(.a(ING186 ), .O(G186));
  buffer g0968(.a(ING189 ), .O(G189));
  buffer g0969(.a(ING190 ), .O(G190));
  buffer g0970(.a(ING191 ), .O(G191));
  buffer g0971(.a(ING192 ), .O(G192));
  buffer g0972(.a(ING193 ), .O(G193));
  buffer g0973(.a(ING194 ), .O(G194));
  buffer g0974(.a(ING195 ), .O(G195));
  buffer g0975(.a(ING196 ), .O(G196));
  buffer g0976(.a(ING197 ), .O(G197));
  buffer g0977(.a(ING198 ), .O(G198));
  buffer g0978(.a(ING199 ), .O(G199));
  buffer g0979(.a(ING200 ), .O(G200));
  buffer g0980(.a(ING201 ), .O(G201));
  buffer g0981(.a(ING202 ), .O(G202));
  buffer g0982(.a(ING203 ), .O(G203));
  buffer g0983(.a(ING204 ), .O(G204));
  buffer g0984(.a(ING205 ), .O(G205));
  buffer g0985(.a(ING206 ), .O(G206));
  buffer g0986(.a(ING207 ), .O(G207));
  buffer g0987(.a(ING208 ), .O(G208));
  buffer g0988(.a(ING209 ), .O(G209));
  buffer g0989(.a(ING210 ), .O(G210));
  buffer g0990(.a(ING211 ), .O(G211));
  buffer g0991(.a(ING212 ), .O(G212));
  buffer g0992(.a(ING213 ), .O(G213));
  buffer g0993(.a(ING214 ), .O(G214));
  buffer g0994(.a(ING215 ), .O(G215));
  buffer g0995(.a(ING239 ), .O(G239));
  buffer g0996(.a(ING240 ), .O(G240));
  buffer g0997(.a(ING241 ), .O(G241));
  buffer g0998(.a(ING242 ), .O(G242));
  buffer g0999(.a(ING243 ), .O(G243));
  buffer g1000(.a(ING244 ), .O(G244));
  buffer g1001(.a(ING245 ), .O(G245));
  buffer g1002(.a(ING246 ), .O(G246));
  buffer g1003(.a(ING247 ), .O(G247));
  buffer g1004(.a(ING248 ), .O(G248));
  buffer g1005(.a(ING249 ), .O(G249));
  buffer g1006(.a(ING250 ), .O(G250));
  buffer g1007(.a(ING251 ), .O(G251));
  buffer g1008(.a(ING252 ), .O(G252));
  buffer g1009(.a(ING253 ), .O(G253));
  buffer g1010(.a(ING254 ), .O(G254));
  buffer g1011(.a(ING255 ), .O(G255));
  buffer g1012(.a(ING256 ), .O(G256));
  buffer g1013(.a(ING257 ), .O(G257));
  buffer g1014(.a(ING262 ), .O(G262));
  buffer g1015(.a(ING263 ), .O(G263));
  buffer g1016(.a(ING264 ), .O(G264));
  buffer g1017(.a(ING265 ), .O(G265));
  buffer g1018(.a(ING266 ), .O(G266));
  buffer g1019(.a(ING267 ), .O(G267));
  buffer g1020(.a(ING268 ), .O(G268));
  buffer g1021(.a(ING269 ), .O(G269));
  buffer g1022(.a(ING270 ), .O(G270));
  buffer g1023(.a(ING271 ), .O(G271));
  buffer g1024(.a(ING272 ), .O(G272));
  buffer g1025(.a(ING273 ), .O(G273));
  buffer g1026(.a(ING274 ), .O(G274));
  buffer g1027(.a(ING275 ), .O(G275));
  buffer g1028(.a(ING276 ), .O(G276));
  buffer g1029(.a(ING277 ), .O(G277));
  buffer g1030(.a(ING278 ), .O(G278));
  buffer g1031(.a(ING279 ), .O(G279));
  buffer g1032(.a(G452), .O(G350));
  buffer g1033(.a(G452), .O(G335));
  buffer g1034(.a(G452), .O(G409));
  buffer g1035(.a(G1083), .O(G369));
  buffer g1036(.a(G1083), .O(G367));
  buffer g1037(.a(G2066), .O(G411));
  buffer g1038(.a(G2066), .O(G337));
  buffer g1039(.a(G2066), .O(G384));
  buffer g1040(.a(G452), .O(G391));
  nor2   g1041(.a(n635), .b(n619), .O(G321));
  nor2   g1042(.a(n638), .b(n637), .O(G280));
  inv1   g1043(.a(n648), .O(G323));
  inv1   g1044(.a(n1132), .O(G331));
endmodule


