// Benchmark "c2670_blif" written by ABC on Sun Mar 24 18:39:13 2019

module c2670_blif  ( 
    G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
    G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
    G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
    G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
    G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
    G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
    G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136,
    G137, G138, G139, G140, G141, G142, ING169 , ING174 , ING177 ,
    ING178 , ING179 , ING180 , ING181 , ING182 , ING183 ,
    ING184 , ING185 , ING186 , ING189 , ING190 , ING191 ,
    ING192 , ING193 , ING194 , ING195 , ING196 , ING197 ,
    ING198 , ING199 , ING200 , ING201 , ING202 , ING203 ,
    ING204 , ING205 , ING206 , ING207 , ING208 , ING209 ,
    ING210 , ING211 , ING212 , ING213 , ING214 , ING215 ,
    ING239 , ING240 , ING241 , ING242 , ING243 , ING244 ,
    ING245 , ING246 , ING247 , ING248 , ING249 , ING250 ,
    ING251 , ING252 , ING253 , ING254 , ING255 , ING256 ,
    ING257 , ING262 , ING263 , ING264 , ING265 , ING266 ,
    ING267 , ING268 , ING269 , ING270 , ING271 , ING272 ,
    ING273 , ING274 , ING275 , ING276 , ING277 , ING278 ,
    ING279 , G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083,
    G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986,
    G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100,
    G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451,
    G2454, G2474, G2678,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G350, G335, G409, G369, G367, G411, G337, G384,
    G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173,
    G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171,
    G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
    G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145,
    G395, G295, G331, G397, G329, G231, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20,
    G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36,
    G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74,
    G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90,
    G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105,
    G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
    G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135,
    G136, G137, G138, G139, G140, G141, G142, ING169 , ING174 ,
    ING177 , ING178 , ING179 , ING180 , ING181 , ING182 ,
    ING183 , ING184 , ING185 , ING186 , ING189 , ING190 ,
    ING191 , ING192 , ING193 , ING194 , ING195 , ING196 ,
    ING197 , ING198 , ING199 , ING200 , ING201 , ING202 ,
    ING203 , ING204 , ING205 , ING206 , ING207 , ING208 ,
    ING209 , ING210 , ING211 , ING212 , ING213 , ING214 ,
    ING215 , ING239 , ING240 , ING241 , ING242 , ING243 ,
    ING244 , ING245 , ING246 , ING247 , ING248 , ING249 ,
    ING250 , ING251 , ING252 , ING253 , ING254 , ING255 ,
    ING256 , ING257 , ING262 , ING263 , ING264 , ING265 ,
    ING266 , ING267 , ING268 , ING269 , ING270 , ING271 ,
    ING272 , ING273 , ING274 , ING275 , ING276 , ING277 ,
    ING278 , ING279 , G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185,
    G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199,
    G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211,
    G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
    G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262,
    G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274,
    G275, G276, G277, G278, G279, G350, G335, G409, G369, G367, G411, G337,
    G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391,
    G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168,
    G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284,
    G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
    G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire n382, n383, n384, n385, n386, n387, n388, n389, n390, n392, n393,
    n394, n395, n396, n397, n399, n400, n402, n403, n405, n406, n408, n409,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n425, n426, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
    n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n476, n477,
    n478, n479, n480, n481, n482, n483, n484, n485, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n513, n514, n515, n516,
    n517, n518, n519, n520, n522, n523, n524, n525, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n553, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n565, n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n593, n594, n595, n597, n598, n599,
    n600, n602, n603, n604, n605, n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n626,
    n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
    n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n674, n675,
    n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
    n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
    n700, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743, n744, n745, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n971, n972, n973, n974, n975, n976, n977, n978, n979,
    n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
    n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257;
  inv1   g000(.a(G44), .O(G218));
  inv1   g001(.a(G132), .O(G219));
  inv1   g002(.a(G82), .O(G220));
  inv1   g003(.a(G96), .O(G221));
  inv1   g004(.a(G69), .O(G235));
  inv1   g005(.a(G120), .O(G236));
  inv1   g006(.a(G57), .O(G237));
  inv1   g007(.a(G108), .O(G238));
  inv1   g008(.a(G2072), .O(n382));
  inv1   g009(.a(G2078), .O(n383));
  nor2   g010(.a(n383), .b(n382), .O(n384));
  inv1   g011(.a(n384), .O(n385));
  inv1   g012(.a(G2084), .O(n386));
  inv1   g013(.a(G2090), .O(n387));
  nor2   g014(.a(n387), .b(n386), .O(n388));
  inv1   g015(.a(n388), .O(n389));
  nor2   g016(.a(n389), .b(n385), .O(n390));
  inv1   g017(.a(n390), .O(G158));
  inv1   g018(.a(G661), .O(n392));
  inv1   g019(.a(G2), .O(n393));
  inv1   g020(.a(G15), .O(n394));
  nor2   g021(.a(n394), .b(n393), .O(n395));
  inv1   g022(.a(n395), .O(n396));
  nor2   g023(.a(n396), .b(n392), .O(n397));
  inv1   g024(.a(n397), .O(G259));
  inv1   g025(.a(G94), .O(n399));
  inv1   g026(.a(G452), .O(n400));
  nor2   g027(.a(n400), .b(n399), .O(G173));
  inv1   g028(.a(G7), .O(n402));
  nor2   g029(.a(n392), .b(n402), .O(n403));
  inv1   g030(.a(n403), .O(G223));
  inv1   g031(.a(G567), .O(n405));
  nor2   g032(.a(G223), .b(n405), .O(n406));
  inv1   g033(.a(n406), .O(G234));
  inv1   g034(.a(G2106), .O(n408));
  nor2   g035(.a(G223), .b(n408), .O(n409));
  inv1   g036(.a(n409), .O(G217));
  nor2   g037(.a(G235), .b(G237), .O(n411));
  inv1   g038(.a(n411), .O(n412));
  nor2   g039(.a(G236), .b(G238), .O(n413));
  inv1   g040(.a(n413), .O(n414));
  nor2   g041(.a(n414), .b(n412), .O(n415));
  inv1   g042(.a(n415), .O(n416));
  nor2   g043(.a(G220), .b(G218), .O(n417));
  inv1   g044(.a(n417), .O(n418));
  nor2   g045(.a(G219), .b(G221), .O(n419));
  inv1   g046(.a(n419), .O(n420));
  nor2   g047(.a(n420), .b(n418), .O(n421));
  inv1   g048(.a(n421), .O(n422));
  nor2   g049(.a(n422), .b(n416), .O(G325));
  inv1   g050(.a(G325), .O(G261));
  nor2   g051(.a(n421), .b(n408), .O(n425));
  nor2   g052(.a(n415), .b(n405), .O(n426));
  nor2   g053(.a(n426), .b(n425), .O(G319));
  inv1   g054(.a(G2104), .O(n428));
  nor2   g055(.a(n428), .b(G113), .O(n429));
  inv1   g056(.a(G2105), .O(n430));
  nor2   g057(.a(G2104), .b(G125), .O(n431));
  nor2   g058(.a(n431), .b(n430), .O(n432));
  inv1   g059(.a(n432), .O(n433));
  nor2   g060(.a(n433), .b(n429), .O(n434));
  nor2   g061(.a(n428), .b(G101), .O(n435));
  nor2   g062(.a(G2104), .b(G137), .O(n436));
  nor2   g063(.a(n436), .b(G2105), .O(n437));
  inv1   g064(.a(n437), .O(n438));
  nor2   g065(.a(n438), .b(n435), .O(n439));
  nor2   g066(.a(n439), .b(n434), .O(G160));
  nor2   g067(.a(n428), .b(G112), .O(n441));
  nor2   g068(.a(G2104), .b(G124), .O(n442));
  nor2   g069(.a(n442), .b(n430), .O(n443));
  inv1   g070(.a(n443), .O(n444));
  nor2   g071(.a(n444), .b(n441), .O(n445));
  nor2   g072(.a(n428), .b(G100), .O(n446));
  nor2   g073(.a(G2104), .b(G136), .O(n447));
  nor2   g074(.a(n447), .b(G2105), .O(n448));
  inv1   g075(.a(n448), .O(n449));
  nor2   g076(.a(n449), .b(n446), .O(n450));
  nor2   g077(.a(n450), .b(n445), .O(G162));
  nor2   g078(.a(n428), .b(G114), .O(n452));
  nor2   g079(.a(G2104), .b(G126), .O(n453));
  nor2   g080(.a(n453), .b(n430), .O(n454));
  inv1   g081(.a(n454), .O(n455));
  nor2   g082(.a(n455), .b(n452), .O(n456));
  nor2   g083(.a(n428), .b(G102), .O(n457));
  nor2   g084(.a(G2104), .b(G138), .O(n458));
  nor2   g085(.a(n458), .b(G2105), .O(n459));
  inv1   g086(.a(n459), .O(n460));
  nor2   g087(.a(n460), .b(n457), .O(n461));
  nor2   g088(.a(n461), .b(n456), .O(G164));
  inv1   g089(.a(G543), .O(n463));
  nor2   g090(.a(n463), .b(G75), .O(n464));
  inv1   g091(.a(G651), .O(n465));
  nor2   g092(.a(G543), .b(G62), .O(n466));
  nor2   g093(.a(n466), .b(n465), .O(n467));
  inv1   g094(.a(n467), .O(n468));
  nor2   g095(.a(n468), .b(n464), .O(n469));
  nor2   g096(.a(n463), .b(G50), .O(n470));
  nor2   g097(.a(G543), .b(G88), .O(n471));
  nor2   g098(.a(n471), .b(G651), .O(n472));
  inv1   g099(.a(n472), .O(n473));
  nor2   g100(.a(n473), .b(n470), .O(n474));
  nor2   g101(.a(n474), .b(n469), .O(G166));
  nor2   g102(.a(n463), .b(G76), .O(n476));
  nor2   g103(.a(G543), .b(G63), .O(n477));
  nor2   g104(.a(n477), .b(n465), .O(n478));
  inv1   g105(.a(n478), .O(n479));
  nor2   g106(.a(n479), .b(n476), .O(n480));
  nor2   g107(.a(n463), .b(G51), .O(n481));
  nor2   g108(.a(G543), .b(G89), .O(n482));
  nor2   g109(.a(n482), .b(G651), .O(n483));
  inv1   g110(.a(n483), .O(n484));
  nor2   g111(.a(n484), .b(n481), .O(n485));
  nor2   g112(.a(n485), .b(n480), .O(G168));
  nor2   g113(.a(n463), .b(G77), .O(n487));
  nor2   g114(.a(G543), .b(G64), .O(n488));
  nor2   g115(.a(n488), .b(n465), .O(n489));
  inv1   g116(.a(n489), .O(n490));
  nor2   g117(.a(n490), .b(n487), .O(n491));
  nor2   g118(.a(n463), .b(G52), .O(n492));
  nor2   g119(.a(G543), .b(G90), .O(n493));
  nor2   g120(.a(n493), .b(G651), .O(n494));
  inv1   g121(.a(n494), .O(n495));
  nor2   g122(.a(n495), .b(n492), .O(n496));
  nor2   g123(.a(n496), .b(n491), .O(G171));
  inv1   g124(.a(G860), .O(n498));
  nor2   g125(.a(n463), .b(G68), .O(n499));
  nor2   g126(.a(G543), .b(G56), .O(n500));
  nor2   g127(.a(n500), .b(n465), .O(n501));
  inv1   g128(.a(n501), .O(n502));
  nor2   g129(.a(n502), .b(n499), .O(n503));
  nor2   g130(.a(n463), .b(G43), .O(n504));
  nor2   g131(.a(G543), .b(G81), .O(n505));
  nor2   g132(.a(n505), .b(G651), .O(n506));
  inv1   g133(.a(n506), .O(n507));
  nor2   g134(.a(n507), .b(n504), .O(n508));
  nor2   g135(.a(n508), .b(n503), .O(n509));
  inv1   g136(.a(n509), .O(n510));
  nor2   g137(.a(n510), .b(n498), .O(n511));
  inv1   g138(.a(n511), .O(G153));
  inv1   g139(.a(G36), .O(n513));
  inv1   g140(.a(G319), .O(n514));
  inv1   g141(.a(G483), .O(n515));
  nor2   g142(.a(n392), .b(n515), .O(n516));
  inv1   g143(.a(n516), .O(n517));
  nor2   g144(.a(n517), .b(n514), .O(n518));
  inv1   g145(.a(n518), .O(n519));
  nor2   g146(.a(n519), .b(n513), .O(n520));
  inv1   g147(.a(n520), .O(G176));
  inv1   g148(.a(G1), .O(n522));
  inv1   g149(.a(G3), .O(n523));
  nor2   g150(.a(n523), .b(n522), .O(n524));
  nor2   g151(.a(n524), .b(n519), .O(n525));
  inv1   g152(.a(n525), .O(G188));
  nor2   g153(.a(n463), .b(G78), .O(n527));
  nor2   g154(.a(G543), .b(G65), .O(n528));
  nor2   g155(.a(n528), .b(n465), .O(n529));
  inv1   g156(.a(n529), .O(n530));
  nor2   g157(.a(n530), .b(n527), .O(n531));
  nor2   g158(.a(n463), .b(G53), .O(n532));
  nor2   g159(.a(G543), .b(G91), .O(n533));
  nor2   g160(.a(n533), .b(G651), .O(n534));
  inv1   g161(.a(n534), .O(n535));
  nor2   g162(.a(n535), .b(n532), .O(n536));
  nor2   g163(.a(n536), .b(n531), .O(n537));
  inv1   g164(.a(n537), .O(G299));
  inv1   g165(.a(G171), .O(G301));
  inv1   g166(.a(G168), .O(G286));
  inv1   g167(.a(G166), .O(G303));
  inv1   g168(.a(G74), .O(n542));
  nor2   g169(.a(n465), .b(n542), .O(n543));
  inv1   g170(.a(G49), .O(n544));
  nor2   g171(.a(G651), .b(n544), .O(n545));
  nor2   g172(.a(n545), .b(n463), .O(n546));
  inv1   g173(.a(n546), .O(n547));
  nor2   g174(.a(n547), .b(n543), .O(n548));
  nor2   g175(.a(G543), .b(G87), .O(n549));
  inv1   g176(.a(n549), .O(n550));
  nor2   g177(.a(n550), .b(G651), .O(n551));
  nor2   g178(.a(n551), .b(n548), .O(G288));
  nor2   g179(.a(n463), .b(G73), .O(n553));
  nor2   g180(.a(G543), .b(G61), .O(n554));
  nor2   g181(.a(n554), .b(n465), .O(n555));
  inv1   g182(.a(n555), .O(n556));
  nor2   g183(.a(n556), .b(n553), .O(n557));
  nor2   g184(.a(n463), .b(G48), .O(n558));
  nor2   g185(.a(G543), .b(G86), .O(n559));
  nor2   g186(.a(n559), .b(G651), .O(n560));
  inv1   g187(.a(n560), .O(n561));
  nor2   g188(.a(n561), .b(n558), .O(n562));
  nor2   g189(.a(n562), .b(n557), .O(n563));
  inv1   g190(.a(n563), .O(G305));
  nor2   g191(.a(n463), .b(G72), .O(n565));
  nor2   g192(.a(G543), .b(G60), .O(n566));
  nor2   g193(.a(n566), .b(n465), .O(n567));
  inv1   g194(.a(n567), .O(n568));
  nor2   g195(.a(n568), .b(n565), .O(n569));
  nor2   g196(.a(n463), .b(G47), .O(n570));
  nor2   g197(.a(G543), .b(G85), .O(n571));
  nor2   g198(.a(n571), .b(G651), .O(n572));
  inv1   g199(.a(n572), .O(n573));
  nor2   g200(.a(n573), .b(n570), .O(n574));
  nor2   g201(.a(n574), .b(n569), .O(n575));
  inv1   g202(.a(n575), .O(G290));
  nor2   g203(.a(n463), .b(G79), .O(n577));
  nor2   g204(.a(G543), .b(G66), .O(n578));
  nor2   g205(.a(n578), .b(n465), .O(n579));
  inv1   g206(.a(n579), .O(n580));
  nor2   g207(.a(n580), .b(n577), .O(n581));
  nor2   g208(.a(n463), .b(G54), .O(n582));
  nor2   g209(.a(G543), .b(G92), .O(n583));
  nor2   g210(.a(n583), .b(G651), .O(n584));
  inv1   g211(.a(n584), .O(n585));
  nor2   g212(.a(n585), .b(n582), .O(n586));
  nor2   g213(.a(n586), .b(n581), .O(n587));
  nor2   g214(.a(n587), .b(G868), .O(n588));
  inv1   g215(.a(G868), .O(n589));
  nor2   g216(.a(G171), .b(n589), .O(n590));
  nor2   g217(.a(n590), .b(n588), .O(n591));
  inv1   g218(.a(n591), .O(G284));
  nor2   g219(.a(n537), .b(G868), .O(n593));
  nor2   g220(.a(G168), .b(n589), .O(n594));
  nor2   g221(.a(n594), .b(n593), .O(n595));
  inv1   g222(.a(n595), .O(G297));
  inv1   g223(.a(n587), .O(n597));
  inv1   g224(.a(G559), .O(n598));
  nor2   g225(.a(G860), .b(n598), .O(n599));
  nor2   g226(.a(n599), .b(n597), .O(n600));
  inv1   g227(.a(n600), .O(G148));
  nor2   g228(.a(n597), .b(G559), .O(n602));
  nor2   g229(.a(n602), .b(n589), .O(n603));
  nor2   g230(.a(n509), .b(G868), .O(n604));
  nor2   g231(.a(n604), .b(n603), .O(n605));
  inv1   g232(.a(n605), .O(G282));
  nor2   g233(.a(n428), .b(G111), .O(n607));
  nor2   g234(.a(G2104), .b(G123), .O(n608));
  nor2   g235(.a(n608), .b(n430), .O(n609));
  inv1   g236(.a(n609), .O(n610));
  nor2   g237(.a(n610), .b(n607), .O(n611));
  nor2   g238(.a(n428), .b(G99), .O(n612));
  nor2   g239(.a(G2104), .b(G135), .O(n613));
  nor2   g240(.a(n613), .b(G2105), .O(n614));
  inv1   g241(.a(n614), .O(n615));
  nor2   g242(.a(n615), .b(n612), .O(n616));
  nor2   g243(.a(n616), .b(n611), .O(n617));
  inv1   g244(.a(n617), .O(n618));
  nor2   g245(.a(n618), .b(G2096), .O(n619));
  inv1   g246(.a(G2096), .O(n620));
  nor2   g247(.a(n617), .b(n620), .O(n621));
  nor2   g248(.a(n621), .b(G2100), .O(n622));
  inv1   g249(.a(n622), .O(n623));
  nor2   g250(.a(n623), .b(n619), .O(n624));
  inv1   g251(.a(n624), .O(G156));
  inv1   g252(.a(G2451), .O(n626));
  nor2   g253(.a(G2454), .b(n626), .O(n627));
  inv1   g254(.a(G2454), .O(n628));
  nor2   g255(.a(n628), .b(G2451), .O(n629));
  nor2   g256(.a(n629), .b(n627), .O(n630));
  inv1   g257(.a(n630), .O(n631));
  inv1   g258(.a(G1341), .O(n632));
  nor2   g259(.a(G2427), .b(n632), .O(n633));
  inv1   g260(.a(G2427), .O(n634));
  nor2   g261(.a(n634), .b(G1341), .O(n635));
  nor2   g262(.a(n635), .b(n633), .O(n636));
  inv1   g263(.a(n636), .O(n637));
  nor2   g264(.a(n637), .b(n631), .O(n638));
  nor2   g265(.a(n636), .b(n630), .O(n639));
  nor2   g266(.a(n639), .b(n638), .O(n640));
  inv1   g267(.a(G2443), .O(n641));
  nor2   g268(.a(G2446), .b(n641), .O(n642));
  inv1   g269(.a(G2446), .O(n643));
  nor2   g270(.a(n643), .b(G2443), .O(n644));
  nor2   g271(.a(n644), .b(n642), .O(n645));
  inv1   g272(.a(n645), .O(n646));
  inv1   g273(.a(G1348), .O(n647));
  nor2   g274(.a(G2430), .b(n647), .O(n648));
  inv1   g275(.a(G2430), .O(n649));
  nor2   g276(.a(n649), .b(G1348), .O(n650));
  nor2   g277(.a(n650), .b(n648), .O(n651));
  inv1   g278(.a(n651), .O(n652));
  nor2   g279(.a(G2438), .b(G2435), .O(n653));
  inv1   g280(.a(G2435), .O(n654));
  inv1   g281(.a(G2438), .O(n655));
  nor2   g282(.a(n655), .b(n654), .O(n656));
  nor2   g283(.a(n656), .b(n653), .O(n657));
  nor2   g284(.a(n657), .b(n652), .O(n658));
  inv1   g285(.a(n657), .O(n659));
  nor2   g286(.a(n659), .b(n651), .O(n660));
  nor2   g287(.a(n660), .b(n658), .O(n661));
  inv1   g288(.a(n661), .O(n662));
  nor2   g289(.a(n662), .b(n646), .O(n663));
  nor2   g290(.a(n661), .b(n645), .O(n664));
  nor2   g291(.a(n664), .b(n663), .O(n665));
  nor2   g292(.a(n665), .b(n640), .O(n666));
  inv1   g293(.a(G14), .O(n667));
  inv1   g294(.a(n640), .O(n668));
  inv1   g295(.a(n665), .O(n669));
  nor2   g296(.a(n669), .b(n668), .O(n670));
  nor2   g297(.a(n670), .b(n667), .O(n671));
  inv1   g298(.a(n671), .O(n672));
  nor2   g299(.a(n672), .b(n666), .O(G401));
  inv1   g300(.a(G2678), .O(n674));
  inv1   g301(.a(G2067), .O(n675));
  nor2   g302(.a(G2100), .b(n620), .O(n676));
  inv1   g303(.a(G2100), .O(n677));
  nor2   g304(.a(n677), .b(G2096), .O(n678));
  nor2   g305(.a(n678), .b(n676), .O(n679));
  inv1   g306(.a(n679), .O(n680));
  nor2   g307(.a(n680), .b(n675), .O(n681));
  nor2   g308(.a(n679), .b(G2067), .O(n682));
  nor2   g309(.a(n682), .b(n681), .O(n683));
  nor2   g310(.a(n683), .b(n674), .O(n684));
  inv1   g311(.a(n683), .O(n685));
  nor2   g312(.a(n685), .b(G2678), .O(n686));
  nor2   g313(.a(n686), .b(n684), .O(n687));
  inv1   g314(.a(n687), .O(n688));
  nor2   g315(.a(G2090), .b(G2084), .O(n689));
  nor2   g316(.a(n689), .b(n388), .O(n690));
  inv1   g317(.a(n690), .O(n691));
  nor2   g318(.a(G2078), .b(G2072), .O(n692));
  nor2   g319(.a(n692), .b(n384), .O(n693));
  nor2   g320(.a(n693), .b(n691), .O(n694));
  inv1   g321(.a(n693), .O(n695));
  nor2   g322(.a(n695), .b(n690), .O(n696));
  nor2   g323(.a(n696), .b(n694), .O(n697));
  inv1   g324(.a(n697), .O(n698));
  nor2   g325(.a(n698), .b(n688), .O(n699));
  nor2   g326(.a(n697), .b(n687), .O(n700));
  nor2   g327(.a(n700), .b(n699), .O(G227));
  inv1   g328(.a(G1971), .O(n702));
  nor2   g329(.a(G1976), .b(n702), .O(n703));
  inv1   g330(.a(G1976), .O(n704));
  nor2   g331(.a(n704), .b(G1971), .O(n705));
  nor2   g332(.a(n705), .b(n703), .O(n706));
  inv1   g333(.a(n706), .O(n707));
  inv1   g334(.a(G1991), .O(n708));
  inv1   g335(.a(G1961), .O(n709));
  nor2   g336(.a(G1966), .b(n709), .O(n710));
  inv1   g337(.a(G1966), .O(n711));
  nor2   g338(.a(n711), .b(G1961), .O(n712));
  nor2   g339(.a(n712), .b(n710), .O(n713));
  inv1   g340(.a(n713), .O(n714));
  nor2   g341(.a(n714), .b(n708), .O(n715));
  nor2   g342(.a(n713), .b(G1991), .O(n716));
  nor2   g343(.a(n716), .b(n715), .O(n717));
  nor2   g344(.a(n717), .b(n707), .O(n718));
  inv1   g345(.a(n717), .O(n719));
  nor2   g346(.a(n719), .b(n706), .O(n720));
  nor2   g347(.a(n720), .b(n718), .O(n721));
  inv1   g348(.a(n721), .O(n722));
  inv1   g349(.a(G2474), .O(n723));
  nor2   g350(.a(G1996), .b(G1956), .O(n724));
  inv1   g351(.a(G1956), .O(n725));
  inv1   g352(.a(G1996), .O(n726));
  nor2   g353(.a(n726), .b(n725), .O(n727));
  nor2   g354(.a(n727), .b(n724), .O(n728));
  inv1   g355(.a(n728), .O(n729));
  nor2   g356(.a(n729), .b(n723), .O(n730));
  nor2   g357(.a(n728), .b(G2474), .O(n731));
  nor2   g358(.a(n731), .b(n730), .O(n732));
  inv1   g359(.a(n732), .O(n733));
  inv1   g360(.a(G1981), .O(n734));
  nor2   g361(.a(G1986), .b(n734), .O(n735));
  inv1   g362(.a(G1986), .O(n736));
  nor2   g363(.a(n736), .b(G1981), .O(n737));
  nor2   g364(.a(n737), .b(n735), .O(n738));
  nor2   g365(.a(n738), .b(n733), .O(n739));
  inv1   g366(.a(n738), .O(n740));
  nor2   g367(.a(n740), .b(n732), .O(n741));
  nor2   g368(.a(n741), .b(n739), .O(n742));
  inv1   g369(.a(n742), .O(n743));
  nor2   g370(.a(n743), .b(n722), .O(n744));
  nor2   g371(.a(n742), .b(n721), .O(n745));
  nor2   g372(.a(n745), .b(n744), .O(G229));
  inv1   g373(.a(G6), .O(n747));
  nor2   g374(.a(G16), .b(n747), .O(n748));
  inv1   g375(.a(G16), .O(n749));
  nor2   g376(.a(n563), .b(n749), .O(n750));
  nor2   g377(.a(n750), .b(n748), .O(n751));
  nor2   g378(.a(n751), .b(n734), .O(n752));
  inv1   g379(.a(G26), .O(n753));
  nor2   g380(.a(G29), .b(n753), .O(n754));
  inv1   g381(.a(G29), .O(n755));
  nor2   g382(.a(n428), .b(G116), .O(n756));
  nor2   g383(.a(G2104), .b(G128), .O(n757));
  nor2   g384(.a(n757), .b(n430), .O(n758));
  inv1   g385(.a(n758), .O(n759));
  nor2   g386(.a(n759), .b(n756), .O(n760));
  nor2   g387(.a(n428), .b(G104), .O(n761));
  nor2   g388(.a(G2104), .b(G140), .O(n762));
  nor2   g389(.a(n762), .b(G2105), .O(n763));
  inv1   g390(.a(n763), .O(n764));
  nor2   g391(.a(n764), .b(n761), .O(n765));
  nor2   g392(.a(n765), .b(n760), .O(n766));
  nor2   g393(.a(n766), .b(n755), .O(n767));
  nor2   g394(.a(n767), .b(n754), .O(n768));
  inv1   g395(.a(n768), .O(n769));
  nor2   g396(.a(n769), .b(G2067), .O(n770));
  nor2   g397(.a(n768), .b(n675), .O(n771));
  nor2   g398(.a(n771), .b(n770), .O(n772));
  inv1   g399(.a(n772), .O(n773));
  nor2   g400(.a(n773), .b(n752), .O(n774));
  inv1   g401(.a(n774), .O(n775));
  inv1   g402(.a(G34), .O(n776));
  nor2   g403(.a(n776), .b(G29), .O(n777));
  nor2   g404(.a(G160), .b(n755), .O(n778));
  nor2   g405(.a(n778), .b(n777), .O(n779));
  inv1   g406(.a(n779), .O(n780));
  nor2   g407(.a(n780), .b(G2084), .O(n781));
  inv1   g408(.a(G19), .O(n782));
  nor2   g409(.a(n782), .b(G16), .O(n783));
  nor2   g410(.a(n509), .b(n749), .O(n784));
  nor2   g411(.a(n784), .b(n783), .O(n785));
  inv1   g412(.a(n785), .O(n786));
  nor2   g413(.a(n786), .b(G1341), .O(n787));
  nor2   g414(.a(n787), .b(n781), .O(n788));
  inv1   g415(.a(n788), .O(n789));
  inv1   g416(.a(G35), .O(n790));
  nor2   g417(.a(n790), .b(G29), .O(n791));
  nor2   g418(.a(G162), .b(n755), .O(n792));
  nor2   g419(.a(n792), .b(n791), .O(n793));
  nor2   g420(.a(n793), .b(n387), .O(n794));
  nor2   g421(.a(n785), .b(n632), .O(n795));
  nor2   g422(.a(n795), .b(n794), .O(n796));
  inv1   g423(.a(n796), .O(n797));
  nor2   g424(.a(n797), .b(n789), .O(n798));
  inv1   g425(.a(n798), .O(n799));
  inv1   g426(.a(n793), .O(n800));
  nor2   g427(.a(n800), .b(G2090), .O(n801));
  inv1   g428(.a(G21), .O(n802));
  nor2   g429(.a(n802), .b(G16), .O(n803));
  nor2   g430(.a(G168), .b(n749), .O(n804));
  nor2   g431(.a(n804), .b(n803), .O(n805));
  nor2   g432(.a(n805), .b(n711), .O(n806));
  nor2   g433(.a(n806), .b(n801), .O(n807));
  inv1   g434(.a(n807), .O(n808));
  inv1   g435(.a(G25), .O(n809));
  nor2   g436(.a(G29), .b(n809), .O(n810));
  nor2   g437(.a(n428), .b(G107), .O(n811));
  nor2   g438(.a(G2104), .b(G119), .O(n812));
  nor2   g439(.a(n812), .b(n430), .O(n813));
  inv1   g440(.a(n813), .O(n814));
  nor2   g441(.a(n814), .b(n811), .O(n815));
  nor2   g442(.a(n428), .b(G95), .O(n816));
  nor2   g443(.a(G2104), .b(G131), .O(n817));
  nor2   g444(.a(n817), .b(G2105), .O(n818));
  inv1   g445(.a(n818), .O(n819));
  nor2   g446(.a(n819), .b(n816), .O(n820));
  nor2   g447(.a(n820), .b(n815), .O(n821));
  nor2   g448(.a(n821), .b(n755), .O(n822));
  nor2   g449(.a(n822), .b(n810), .O(n823));
  inv1   g450(.a(n823), .O(n824));
  nor2   g451(.a(n824), .b(G1991), .O(n825));
  nor2   g452(.a(n823), .b(n708), .O(n826));
  nor2   g453(.a(n826), .b(n825), .O(n827));
  inv1   g454(.a(n827), .O(n828));
  nor2   g455(.a(n828), .b(n808), .O(n829));
  inv1   g456(.a(n829), .O(n830));
  nor2   g457(.a(n830), .b(n799), .O(n831));
  inv1   g458(.a(n831), .O(n832));
  nor2   g459(.a(n832), .b(n775), .O(n833));
  inv1   g460(.a(n833), .O(n834));
  nor2   g461(.a(G288), .b(n749), .O(n835));
  nor2   g462(.a(G23), .b(G16), .O(n836));
  nor2   g463(.a(n836), .b(n835), .O(n837));
  nor2   g464(.a(n837), .b(n704), .O(n838));
  inv1   g465(.a(n837), .O(n839));
  nor2   g466(.a(n839), .b(G1976), .O(n840));
  nor2   g467(.a(n840), .b(n838), .O(n841));
  inv1   g468(.a(G20), .O(n842));
  nor2   g469(.a(n842), .b(G16), .O(n843));
  nor2   g470(.a(n537), .b(n749), .O(n844));
  nor2   g471(.a(n844), .b(n843), .O(n845));
  nor2   g472(.a(n845), .b(G1956), .O(n846));
  inv1   g473(.a(n845), .O(n847));
  nor2   g474(.a(n847), .b(n725), .O(n848));
  nor2   g475(.a(n848), .b(n846), .O(n849));
  inv1   g476(.a(G32), .O(n850));
  nor2   g477(.a(n850), .b(G29), .O(n851));
  nor2   g478(.a(n428), .b(G117), .O(n852));
  nor2   g479(.a(G2104), .b(G129), .O(n853));
  nor2   g480(.a(n853), .b(n430), .O(n854));
  inv1   g481(.a(n854), .O(n855));
  nor2   g482(.a(n855), .b(n852), .O(n856));
  nor2   g483(.a(n428), .b(G105), .O(n857));
  nor2   g484(.a(G2104), .b(G141), .O(n858));
  nor2   g485(.a(n858), .b(G2105), .O(n859));
  inv1   g486(.a(n859), .O(n860));
  nor2   g487(.a(n860), .b(n857), .O(n861));
  nor2   g488(.a(n861), .b(n856), .O(n862));
  nor2   g489(.a(n862), .b(n755), .O(n863));
  nor2   g490(.a(n863), .b(n851), .O(n864));
  nor2   g491(.a(n864), .b(G1996), .O(n865));
  inv1   g492(.a(n864), .O(n866));
  nor2   g493(.a(n866), .b(n726), .O(n867));
  nor2   g494(.a(n867), .b(n865), .O(n868));
  nor2   g495(.a(n868), .b(n849), .O(n869));
  inv1   g496(.a(n869), .O(n870));
  nor2   g497(.a(n870), .b(n841), .O(n871));
  inv1   g498(.a(n871), .O(n872));
  inv1   g499(.a(n751), .O(n873));
  nor2   g500(.a(n873), .b(G1981), .O(n874));
  inv1   g501(.a(G27), .O(n875));
  nor2   g502(.a(G29), .b(n875), .O(n876));
  nor2   g503(.a(G164), .b(n755), .O(n877));
  nor2   g504(.a(n877), .b(n876), .O(n878));
  nor2   g505(.a(n878), .b(n383), .O(n879));
  nor2   g506(.a(n879), .b(n874), .O(n880));
  inv1   g507(.a(n880), .O(n881));
  inv1   g508(.a(G24), .O(n882));
  nor2   g509(.a(n882), .b(G16), .O(n883));
  nor2   g510(.a(n575), .b(n749), .O(n884));
  nor2   g511(.a(n884), .b(n883), .O(n885));
  nor2   g512(.a(n885), .b(n736), .O(n886));
  inv1   g513(.a(n885), .O(n887));
  nor2   g514(.a(n887), .b(G1986), .O(n888));
  nor2   g515(.a(n888), .b(n886), .O(n889));
  inv1   g516(.a(n889), .O(n890));
  nor2   g517(.a(n890), .b(n881), .O(n891));
  inv1   g518(.a(n891), .O(n892));
  inv1   g519(.a(G4), .O(n893));
  nor2   g520(.a(G16), .b(n893), .O(n894));
  nor2   g521(.a(n587), .b(n749), .O(n895));
  nor2   g522(.a(n895), .b(n894), .O(n896));
  nor2   g523(.a(n896), .b(G1348), .O(n897));
  inv1   g524(.a(n896), .O(n898));
  nor2   g525(.a(n898), .b(n647), .O(n899));
  nor2   g526(.a(n899), .b(n897), .O(n900));
  inv1   g527(.a(n878), .O(n901));
  nor2   g528(.a(n901), .b(G2078), .O(n902));
  nor2   g529(.a(n618), .b(n755), .O(n903));
  inv1   g530(.a(G11), .O(n904));
  nor2   g531(.a(G29), .b(G28), .O(n905));
  nor2   g532(.a(n905), .b(n904), .O(n906));
  inv1   g533(.a(n906), .O(n907));
  nor2   g534(.a(n907), .b(n903), .O(n908));
  inv1   g535(.a(n908), .O(n909));
  nor2   g536(.a(n909), .b(n902), .O(n910));
  inv1   g537(.a(n910), .O(n911));
  nor2   g538(.a(n911), .b(n900), .O(n912));
  inv1   g539(.a(n912), .O(n913));
  nor2   g540(.a(n913), .b(n892), .O(n914));
  inv1   g541(.a(n914), .O(n915));
  nor2   g542(.a(n779), .b(n386), .O(n916));
  inv1   g543(.a(n805), .O(n917));
  nor2   g544(.a(n917), .b(G1966), .O(n918));
  nor2   g545(.a(n918), .b(n916), .O(n919));
  inv1   g546(.a(n919), .O(n920));
  inv1   g547(.a(G33), .O(n921));
  nor2   g548(.a(n921), .b(G29), .O(n922));
  nor2   g549(.a(n428), .b(G115), .O(n923));
  nor2   g550(.a(G2104), .b(G127), .O(n924));
  nor2   g551(.a(n924), .b(n430), .O(n925));
  inv1   g552(.a(n925), .O(n926));
  nor2   g553(.a(n926), .b(n923), .O(n927));
  nor2   g554(.a(n428), .b(G103), .O(n928));
  nor2   g555(.a(G2104), .b(G139), .O(n929));
  nor2   g556(.a(n929), .b(G2105), .O(n930));
  inv1   g557(.a(n930), .O(n931));
  nor2   g558(.a(n931), .b(n928), .O(n932));
  nor2   g559(.a(n932), .b(n927), .O(n933));
  nor2   g560(.a(n933), .b(n755), .O(n934));
  nor2   g561(.a(n934), .b(n922), .O(n935));
  nor2   g562(.a(n935), .b(n382), .O(n936));
  inv1   g563(.a(n935), .O(n937));
  nor2   g564(.a(n937), .b(G2072), .O(n938));
  nor2   g565(.a(n938), .b(n936), .O(n939));
  inv1   g566(.a(n939), .O(n940));
  nor2   g567(.a(n940), .b(n920), .O(n941));
  inv1   g568(.a(n941), .O(n942));
  inv1   g569(.a(G22), .O(n943));
  nor2   g570(.a(n943), .b(G16), .O(n944));
  nor2   g571(.a(G166), .b(n749), .O(n945));
  nor2   g572(.a(n945), .b(n944), .O(n946));
  nor2   g573(.a(n946), .b(n702), .O(n947));
  inv1   g574(.a(n946), .O(n948));
  nor2   g575(.a(n948), .b(G1971), .O(n949));
  nor2   g576(.a(n949), .b(n947), .O(n950));
  inv1   g577(.a(n950), .O(n951));
  inv1   g578(.a(G5), .O(n952));
  nor2   g579(.a(G16), .b(n952), .O(n953));
  nor2   g580(.a(G171), .b(n749), .O(n954));
  nor2   g581(.a(n954), .b(n953), .O(n955));
  nor2   g582(.a(n955), .b(n709), .O(n956));
  inv1   g583(.a(n955), .O(n957));
  nor2   g584(.a(n957), .b(G1961), .O(n958));
  nor2   g585(.a(n958), .b(n956), .O(n959));
  inv1   g586(.a(n959), .O(n960));
  nor2   g587(.a(n960), .b(n951), .O(n961));
  inv1   g588(.a(n961), .O(n962));
  nor2   g589(.a(n962), .b(n942), .O(n963));
  inv1   g590(.a(n963), .O(n964));
  nor2   g591(.a(n964), .b(n915), .O(n965));
  inv1   g592(.a(n965), .O(n966));
  nor2   g593(.a(n966), .b(n872), .O(n967));
  inv1   g594(.a(n967), .O(n968));
  nor2   g595(.a(n968), .b(n834), .O(G311));
  inv1   g596(.a(G311), .O(G150));
  inv1   g597(.a(n599), .O(n971));
  nor2   g598(.a(n971), .b(n597), .O(n972));
  nor2   g599(.a(n972), .b(n511), .O(n973));
  inv1   g600(.a(n973), .O(n974));
  nor2   g601(.a(n463), .b(G80), .O(n975));
  nor2   g602(.a(G543), .b(G67), .O(n976));
  nor2   g603(.a(n976), .b(n465), .O(n977));
  inv1   g604(.a(n977), .O(n978));
  nor2   g605(.a(n978), .b(n975), .O(n979));
  nor2   g606(.a(n463), .b(G55), .O(n980));
  nor2   g607(.a(G543), .b(G93), .O(n981));
  nor2   g608(.a(n981), .b(G651), .O(n982));
  inv1   g609(.a(n982), .O(n983));
  nor2   g610(.a(n983), .b(n980), .O(n984));
  nor2   g611(.a(n984), .b(n979), .O(n985));
  nor2   g612(.a(n985), .b(n510), .O(n986));
  inv1   g613(.a(n985), .O(n987));
  nor2   g614(.a(n987), .b(n509), .O(n988));
  nor2   g615(.a(n988), .b(n986), .O(n989));
  inv1   g616(.a(n989), .O(n990));
  nor2   g617(.a(n990), .b(n974), .O(n991));
  nor2   g618(.a(n989), .b(n973), .O(n992));
  nor2   g619(.a(n992), .b(n991), .O(n993));
  inv1   g620(.a(n993), .O(G145));
  inv1   g621(.a(G160), .O(n995));
  nor2   g622(.a(G162), .b(n995), .O(n996));
  inv1   g623(.a(G162), .O(n997));
  nor2   g624(.a(n997), .b(G160), .O(n998));
  nor2   g625(.a(n998), .b(n996), .O(n999));
  inv1   g626(.a(n999), .O(n1000));
  nor2   g627(.a(n1000), .b(n618), .O(n1001));
  nor2   g628(.a(n999), .b(n617), .O(n1002));
  nor2   g629(.a(n1002), .b(n1001), .O(n1003));
  inv1   g630(.a(n821), .O(n1004));
  nor2   g631(.a(n428), .b(G118), .O(n1005));
  nor2   g632(.a(G2104), .b(G130), .O(n1006));
  nor2   g633(.a(n1006), .b(n430), .O(n1007));
  inv1   g634(.a(n1007), .O(n1008));
  nor2   g635(.a(n1008), .b(n1005), .O(n1009));
  nor2   g636(.a(n428), .b(G106), .O(n1010));
  nor2   g637(.a(G2104), .b(G142), .O(n1011));
  nor2   g638(.a(n1011), .b(G2105), .O(n1012));
  inv1   g639(.a(n1012), .O(n1013));
  nor2   g640(.a(n1013), .b(n1010), .O(n1014));
  nor2   g641(.a(n1014), .b(n1009), .O(n1015));
  inv1   g642(.a(n1015), .O(n1016));
  nor2   g643(.a(n1016), .b(G164), .O(n1017));
  inv1   g644(.a(G164), .O(n1018));
  nor2   g645(.a(n1015), .b(n1018), .O(n1019));
  nor2   g646(.a(n1019), .b(n1017), .O(n1020));
  nor2   g647(.a(n1020), .b(n1004), .O(n1021));
  inv1   g648(.a(n1020), .O(n1022));
  nor2   g649(.a(n1022), .b(n821), .O(n1023));
  nor2   g650(.a(n1023), .b(n1021), .O(n1024));
  inv1   g651(.a(n1024), .O(n1025));
  inv1   g652(.a(n766), .O(n1026));
  nor2   g653(.a(n933), .b(n862), .O(n1027));
  inv1   g654(.a(n862), .O(n1028));
  inv1   g655(.a(n933), .O(n1029));
  nor2   g656(.a(n1029), .b(n1028), .O(n1030));
  nor2   g657(.a(n1030), .b(n1027), .O(n1031));
  nor2   g658(.a(n1031), .b(n1026), .O(n1032));
  inv1   g659(.a(n1031), .O(n1033));
  nor2   g660(.a(n1033), .b(n766), .O(n1034));
  nor2   g661(.a(n1034), .b(n1032), .O(n1035));
  inv1   g662(.a(n1035), .O(n1036));
  nor2   g663(.a(n1036), .b(n1025), .O(n1037));
  nor2   g664(.a(n1035), .b(n1024), .O(n1038));
  nor2   g665(.a(n1038), .b(n1037), .O(n1039));
  inv1   g666(.a(n1039), .O(n1040));
  nor2   g667(.a(n1040), .b(n1003), .O(n1041));
  inv1   g668(.a(n1003), .O(n1042));
  nor2   g669(.a(n1039), .b(n1042), .O(n1043));
  nor2   g670(.a(n1043), .b(G37), .O(n1044));
  inv1   g671(.a(n1044), .O(n1045));
  nor2   g672(.a(n1045), .b(n1041), .O(G395));
  inv1   g673(.a(n602), .O(n1047));
  nor2   g674(.a(n989), .b(n537), .O(n1048));
  nor2   g675(.a(n990), .b(G299), .O(n1049));
  nor2   g676(.a(n1049), .b(n1048), .O(n1050));
  nor2   g677(.a(n1050), .b(n1047), .O(n1051));
  nor2   g678(.a(n1050), .b(n587), .O(n1052));
  inv1   g679(.a(n1050), .O(n1053));
  nor2   g680(.a(n1053), .b(n597), .O(n1054));
  nor2   g681(.a(n1054), .b(n1052), .O(n1055));
  nor2   g682(.a(n1055), .b(n602), .O(n1056));
  nor2   g683(.a(n1056), .b(n1051), .O(n1057));
  inv1   g684(.a(n1057), .O(n1058));
  nor2   g685(.a(n575), .b(G303), .O(n1059));
  nor2   g686(.a(G290), .b(G166), .O(n1060));
  nor2   g687(.a(n1060), .b(n1059), .O(n1061));
  inv1   g688(.a(n1061), .O(n1062));
  nor2   g689(.a(G305), .b(G288), .O(n1063));
  inv1   g690(.a(G288), .O(n1064));
  nor2   g691(.a(n563), .b(n1064), .O(n1065));
  nor2   g692(.a(n1065), .b(n1063), .O(n1066));
  inv1   g693(.a(n1066), .O(n1067));
  nor2   g694(.a(n1067), .b(n1062), .O(n1068));
  nor2   g695(.a(n1066), .b(n1061), .O(n1069));
  nor2   g696(.a(n1069), .b(n1068), .O(n1070));
  inv1   g697(.a(n1070), .O(n1071));
  nor2   g698(.a(n1071), .b(n1058), .O(n1072));
  nor2   g699(.a(n1070), .b(n1057), .O(n1073));
  nor2   g700(.a(n1073), .b(n1072), .O(n1074));
  nor2   g701(.a(n1074), .b(n589), .O(n1075));
  nor2   g702(.a(n985), .b(G868), .O(n1076));
  nor2   g703(.a(n1076), .b(n1075), .O(n1077));
  inv1   g704(.a(n1077), .O(G295));
  inv1   g705(.a(n1055), .O(n1079));
  nor2   g706(.a(G171), .b(G286), .O(n1080));
  nor2   g707(.a(G301), .b(G168), .O(n1081));
  nor2   g708(.a(n1081), .b(n1080), .O(n1082));
  inv1   g709(.a(n1082), .O(n1083));
  nor2   g710(.a(n1083), .b(n1079), .O(n1084));
  nor2   g711(.a(n1082), .b(n1055), .O(n1085));
  nor2   g712(.a(n1085), .b(n1084), .O(n1086));
  nor2   g713(.a(n1086), .b(n1070), .O(n1087));
  inv1   g714(.a(n1086), .O(n1088));
  nor2   g715(.a(n1088), .b(n1071), .O(n1089));
  nor2   g716(.a(n1089), .b(G37), .O(n1090));
  inv1   g717(.a(n1090), .O(n1091));
  nor2   g718(.a(n1091), .b(n1087), .O(G397));
  nor2   g719(.a(G164), .b(G1384), .O(n1093));
  inv1   g720(.a(n1093), .O(n1094));
  inv1   g721(.a(G40), .O(n1095));
  nor2   g722(.a(n995), .b(n1095), .O(n1096));
  inv1   g723(.a(n1096), .O(n1097));
  nor2   g724(.a(n1097), .b(n1094), .O(n1098));
  nor2   g725(.a(n1098), .b(n711), .O(n1099));
  inv1   g726(.a(G8), .O(n1100));
  inv1   g727(.a(n1098), .O(n1101));
  nor2   g728(.a(n1101), .b(n386), .O(n1102));
  nor2   g729(.a(n1102), .b(n1100), .O(n1103));
  inv1   g730(.a(n1103), .O(n1104));
  nor2   g731(.a(n1104), .b(n1099), .O(n1105));
  nor2   g732(.a(G168), .b(n1100), .O(n1106));
  inv1   g733(.a(n1106), .O(n1107));
  nor2   g734(.a(n1107), .b(n1105), .O(n1108));
  nor2   g735(.a(n1098), .b(n1100), .O(n1109));
  inv1   g736(.a(n1109), .O(n1110));
  nor2   g737(.a(G288), .b(G1976), .O(n1111));
  nor2   g738(.a(n1064), .b(n704), .O(n1112));
  nor2   g739(.a(n563), .b(n734), .O(n1113));
  nor2   g740(.a(n1113), .b(n1112), .O(n1114));
  inv1   g741(.a(n1114), .O(n1115));
  nor2   g742(.a(n1115), .b(n1111), .O(n1116));
  nor2   g743(.a(n1116), .b(n1110), .O(n1117));
  nor2   g744(.a(G305), .b(G1981), .O(n1118));
  inv1   g745(.a(n1118), .O(n1119));
  nor2   g746(.a(n1119), .b(n1110), .O(n1120));
  nor2   g747(.a(n1120), .b(n1117), .O(n1121));
  inv1   g748(.a(n1121), .O(n1122));
  inv1   g749(.a(n1105), .O(n1123));
  nor2   g750(.a(n1123), .b(G286), .O(n1124));
  nor2   g751(.a(n1124), .b(n1122), .O(n1125));
  inv1   g752(.a(n1125), .O(n1126));
  nor2   g753(.a(n1126), .b(n1108), .O(n1127));
  inv1   g754(.a(n1127), .O(n1128));
  nor2   g755(.a(n1098), .b(n702), .O(n1129));
  nor2   g756(.a(n1101), .b(n387), .O(n1130));
  nor2   g757(.a(n1130), .b(n1100), .O(n1131));
  inv1   g758(.a(n1131), .O(n1132));
  nor2   g759(.a(n1132), .b(n1129), .O(n1133));
  nor2   g760(.a(G166), .b(n1100), .O(n1134));
  inv1   g761(.a(n1134), .O(n1135));
  nor2   g762(.a(n1135), .b(n1133), .O(n1136));
  inv1   g763(.a(n1133), .O(n1137));
  nor2   g764(.a(n1137), .b(G303), .O(n1138));
  nor2   g765(.a(n1138), .b(n1136), .O(n1139));
  inv1   g766(.a(n1139), .O(n1140));
  nor2   g767(.a(n1098), .b(n709), .O(n1141));
  nor2   g768(.a(n1101), .b(n383), .O(n1142));
  nor2   g769(.a(n1142), .b(n1141), .O(n1143));
  nor2   g770(.a(n1143), .b(G171), .O(n1144));
  inv1   g771(.a(n1143), .O(n1145));
  nor2   g772(.a(n1145), .b(G301), .O(n1146));
  nor2   g773(.a(n587), .b(n675), .O(n1147));
  nor2   g774(.a(n510), .b(G1996), .O(n1148));
  inv1   g775(.a(n1148), .O(n1149));
  nor2   g776(.a(n1149), .b(n1147), .O(n1150));
  nor2   g777(.a(n597), .b(G2067), .O(n1151));
  nor2   g778(.a(G299), .b(G2072), .O(n1152));
  nor2   g779(.a(n1152), .b(n1151), .O(n1153));
  inv1   g780(.a(n1153), .O(n1154));
  nor2   g781(.a(n1154), .b(n1150), .O(n1155));
  nor2   g782(.a(n537), .b(n382), .O(n1156));
  nor2   g783(.a(n1156), .b(n1101), .O(n1157));
  inv1   g784(.a(n1157), .O(n1158));
  nor2   g785(.a(n1158), .b(n1155), .O(n1159));
  nor2   g786(.a(n587), .b(n647), .O(n1160));
  nor2   g787(.a(n510), .b(G1341), .O(n1161));
  inv1   g788(.a(n1161), .O(n1162));
  nor2   g789(.a(n1162), .b(n1160), .O(n1163));
  nor2   g790(.a(n597), .b(G1348), .O(n1164));
  nor2   g791(.a(G299), .b(G1956), .O(n1165));
  nor2   g792(.a(n1165), .b(n1164), .O(n1166));
  inv1   g793(.a(n1166), .O(n1167));
  nor2   g794(.a(n1167), .b(n1163), .O(n1168));
  nor2   g795(.a(n537), .b(n725), .O(n1169));
  nor2   g796(.a(n1169), .b(n1098), .O(n1170));
  inv1   g797(.a(n1170), .O(n1171));
  nor2   g798(.a(n1171), .b(n1168), .O(n1172));
  nor2   g799(.a(n1172), .b(n1159), .O(n1173));
  nor2   g800(.a(n1173), .b(n1146), .O(n1174));
  inv1   g801(.a(n1174), .O(n1175));
  nor2   g802(.a(n1175), .b(n1144), .O(n1176));
  inv1   g803(.a(n1176), .O(n1177));
  nor2   g804(.a(n1177), .b(n1140), .O(n1178));
  inv1   g805(.a(n1178), .O(n1179));
  nor2   g806(.a(n1179), .b(n1128), .O(n1180));
  inv1   g807(.a(n1146), .O(n1181));
  nor2   g808(.a(n1181), .b(n1140), .O(n1182));
  inv1   g809(.a(n1182), .O(n1183));
  nor2   g810(.a(n1183), .b(n1128), .O(n1184));
  inv1   g811(.a(n1124), .O(n1185));
  nor2   g812(.a(n1185), .b(n1122), .O(n1186));
  inv1   g813(.a(n1186), .O(n1187));
  nor2   g814(.a(n1187), .b(n1140), .O(n1188));
  inv1   g815(.a(n1138), .O(n1189));
  nor2   g816(.a(n1189), .b(n1117), .O(n1190));
  inv1   g817(.a(n1117), .O(n1191));
  nor2   g818(.a(n1191), .b(n1115), .O(n1192));
  nor2   g819(.a(n1192), .b(n1120), .O(n1193));
  inv1   g820(.a(n1193), .O(n1194));
  nor2   g821(.a(n1194), .b(n1190), .O(n1195));
  inv1   g822(.a(n1195), .O(n1196));
  nor2   g823(.a(n1196), .b(n1188), .O(n1197));
  inv1   g824(.a(n1197), .O(n1198));
  nor2   g825(.a(n1198), .b(n1184), .O(n1199));
  inv1   g826(.a(n1199), .O(n1200));
  nor2   g827(.a(n1200), .b(n1180), .O(n1201));
  nor2   g828(.a(n1097), .b(n1093), .O(n1202));
  inv1   g829(.a(n1202), .O(n1203));
  nor2   g830(.a(n1203), .b(G2067), .O(n1204));
  inv1   g831(.a(n1204), .O(n1205));
  nor2   g832(.a(n1205), .b(n1026), .O(n1206));
  nor2   g833(.a(n1204), .b(n766), .O(n1207));
  nor2   g834(.a(n1028), .b(G1996), .O(n1208));
  nor2   g835(.a(n862), .b(n726), .O(n1209));
  nor2   g836(.a(n1209), .b(n1208), .O(n1210));
  inv1   g837(.a(n1210), .O(n1211));
  nor2   g838(.a(n1211), .b(n1207), .O(n1212));
  inv1   g839(.a(n1212), .O(n1213));
  nor2   g840(.a(n1213), .b(n1206), .O(n1214));
  inv1   g841(.a(n1214), .O(n1215));
  nor2   g842(.a(n1203), .b(G1991), .O(n1216));
  inv1   g843(.a(n1216), .O(n1217));
  nor2   g844(.a(n1217), .b(n1004), .O(n1218));
  nor2   g845(.a(n1216), .b(n821), .O(n1219));
  nor2   g846(.a(n1219), .b(n1218), .O(n1220));
  inv1   g847(.a(n1220), .O(n1221));
  nor2   g848(.a(n1221), .b(n1215), .O(n1222));
  inv1   g849(.a(n1222), .O(n1223));
  nor2   g850(.a(G290), .b(G1986), .O(n1224));
  nor2   g851(.a(n575), .b(n736), .O(n1225));
  nor2   g852(.a(n1225), .b(n1224), .O(n1226));
  inv1   g853(.a(n1226), .O(n1227));
  nor2   g854(.a(n1227), .b(n1223), .O(n1228));
  nor2   g855(.a(n1228), .b(n1203), .O(n1229));
  nor2   g856(.a(n1229), .b(n1201), .O(n1230));
  inv1   g857(.a(n1224), .O(n1231));
  nor2   g858(.a(n1231), .b(n1203), .O(n1232));
  inv1   g859(.a(n1232), .O(n1233));
  nor2   g860(.a(n1233), .b(n1223), .O(n1234));
  inv1   g861(.a(n1218), .O(n1235));
  nor2   g862(.a(n1235), .b(n1215), .O(n1236));
  inv1   g863(.a(n1208), .O(n1237));
  nor2   g864(.a(n1237), .b(n1203), .O(n1238));
  inv1   g865(.a(n1238), .O(n1239));
  nor2   g866(.a(n1239), .b(n1207), .O(n1240));
  nor2   g867(.a(n1240), .b(n1206), .O(n1241));
  inv1   g868(.a(n1241), .O(n1242));
  nor2   g869(.a(n1242), .b(n1236), .O(n1243));
  inv1   g870(.a(n1243), .O(n1244));
  nor2   g871(.a(n1244), .b(n1234), .O(n1245));
  inv1   g872(.a(n1245), .O(n1246));
  nor2   g873(.a(n1246), .b(n1230), .O(n1247));
  inv1   g874(.a(n1247), .O(G329));
  nor2   g875(.a(G227), .b(n514), .O(n1250));
  inv1   g876(.a(n1250), .O(n1251));
  nor2   g877(.a(n1251), .b(G229), .O(n1252));
  inv1   g878(.a(n1252), .O(n1253));
  nor2   g879(.a(n1253), .b(G401), .O(n1254));
  inv1   g880(.a(n1254), .O(n1255));
  nor2   g881(.a(n1255), .b(G395), .O(n1256));
  inv1   g882(.a(n1256), .O(n1257));
  nor2   g883(.a(n1257), .b(G397), .O(G308));
  inv1   g884(.a(G308), .O(G225));
  zero   g885(.O(G231));
  buffer g886(.a(ING169 ), .O(G169));
  buffer g887(.a(ING174 ), .O(G174));
  buffer g888(.a(ING177 ), .O(G177));
  buffer g889(.a(ING178 ), .O(G178));
  buffer g890(.a(ING179 ), .O(G179));
  buffer g891(.a(ING180 ), .O(G180));
  buffer g892(.a(ING181 ), .O(G181));
  buffer g893(.a(ING182 ), .O(G182));
  buffer g894(.a(ING183 ), .O(G183));
  buffer g895(.a(ING184 ), .O(G184));
  buffer g896(.a(ING185 ), .O(G185));
  buffer g897(.a(ING186 ), .O(G186));
  buffer g898(.a(ING189 ), .O(G189));
  buffer g899(.a(ING190 ), .O(G190));
  buffer g900(.a(ING191 ), .O(G191));
  buffer g901(.a(ING192 ), .O(G192));
  buffer g902(.a(ING193 ), .O(G193));
  buffer g903(.a(ING194 ), .O(G194));
  buffer g904(.a(ING195 ), .O(G195));
  buffer g905(.a(ING196 ), .O(G196));
  buffer g906(.a(ING197 ), .O(G197));
  buffer g907(.a(ING198 ), .O(G198));
  buffer g908(.a(ING199 ), .O(G199));
  buffer g909(.a(ING200 ), .O(G200));
  buffer g910(.a(ING201 ), .O(G201));
  buffer g911(.a(ING202 ), .O(G202));
  buffer g912(.a(ING203 ), .O(G203));
  buffer g913(.a(ING204 ), .O(G204));
  buffer g914(.a(ING205 ), .O(G205));
  buffer g915(.a(ING206 ), .O(G206));
  buffer g916(.a(ING207 ), .O(G207));
  buffer g917(.a(ING208 ), .O(G208));
  buffer g918(.a(ING209 ), .O(G209));
  buffer g919(.a(ING210 ), .O(G210));
  buffer g920(.a(ING211 ), .O(G211));
  buffer g921(.a(ING212 ), .O(G212));
  buffer g922(.a(ING213 ), .O(G213));
  buffer g923(.a(ING214 ), .O(G214));
  buffer g924(.a(ING215 ), .O(G215));
  buffer g925(.a(ING239 ), .O(G239));
  buffer g926(.a(ING240 ), .O(G240));
  buffer g927(.a(ING241 ), .O(G241));
  buffer g928(.a(ING242 ), .O(G242));
  buffer g929(.a(ING243 ), .O(G243));
  buffer g930(.a(ING244 ), .O(G244));
  buffer g931(.a(ING245 ), .O(G245));
  buffer g932(.a(ING246 ), .O(G246));
  buffer g933(.a(ING247 ), .O(G247));
  buffer g934(.a(ING248 ), .O(G248));
  buffer g935(.a(ING249 ), .O(G249));
  buffer g936(.a(ING250 ), .O(G250));
  buffer g937(.a(ING251 ), .O(G251));
  buffer g938(.a(ING252 ), .O(G252));
  buffer g939(.a(ING253 ), .O(G253));
  buffer g940(.a(ING254 ), .O(G254));
  buffer g941(.a(ING255 ), .O(G255));
  buffer g942(.a(ING256 ), .O(G256));
  buffer g943(.a(ING257 ), .O(G257));
  buffer g944(.a(ING262 ), .O(G262));
  buffer g945(.a(ING263 ), .O(G263));
  buffer g946(.a(ING264 ), .O(G264));
  buffer g947(.a(ING265 ), .O(G265));
  buffer g948(.a(ING266 ), .O(G266));
  buffer g949(.a(ING267 ), .O(G267));
  buffer g950(.a(ING268 ), .O(G268));
  buffer g951(.a(ING269 ), .O(G269));
  buffer g952(.a(ING270 ), .O(G270));
  buffer g953(.a(ING271 ), .O(G271));
  buffer g954(.a(ING272 ), .O(G272));
  buffer g955(.a(ING273 ), .O(G273));
  buffer g956(.a(ING274 ), .O(G274));
  buffer g957(.a(ING275 ), .O(G275));
  buffer g958(.a(ING276 ), .O(G276));
  buffer g959(.a(ING277 ), .O(G277));
  buffer g960(.a(ING278 ), .O(G278));
  buffer g961(.a(ING279 ), .O(G279));
  buffer g962(.a(G452), .O(G350));
  buffer g963(.a(G452), .O(G335));
  buffer g964(.a(G452), .O(G409));
  buffer g965(.a(G1083), .O(G369));
  buffer g966(.a(G1083), .O(G367));
  buffer g967(.a(G2066), .O(G411));
  buffer g968(.a(G2066), .O(G337));
  buffer g969(.a(G2066), .O(G384));
  buffer g970(.a(G452), .O(G391));
  inv1   g971(.a(n591), .O(G321));
  inv1   g972(.a(n595), .O(G280));
  inv1   g973(.a(n605), .O(G323));
  inv1   g974(.a(n1077), .O(G331));
endmodule


