// Benchmark "c499_blif" written by ABC on Sun Apr 14 20:03:44 2019

module c499_blif  ( 
    Gid0, Gid1, Gid2, Gid3, Gid4, Gid5, Gid6, Gid7, Gid8, Gid9, Gid10,
    Gid11, Gid12, Gid13, Gid14, Gid15, Gid16, Gid17, Gid18, Gid19, Gid20,
    Gid21, Gid22, Gid23, Gid24, Gid25, Gid26, Gid27, Gid28, Gid29, Gid30,
    Gid31, Gic0, Gic1, Gic2, Gic3, Gic4, Gic5, Gic6, Gic7, Gr,
    God0, God1, God2, God3, God4, God5, God6, God7, God8, God9, God10,
    God11, God12, God13, God14, God15, God16, God17, God18, God19, God20,
    God21, God22, God23, God24, God25, God26, God27, God28, God29, God30,
    God31  );
  input  Gid0, Gid1, Gid2, Gid3, Gid4, Gid5, Gid6, Gid7, Gid8, Gid9,
    Gid10, Gid11, Gid12, Gid13, Gid14, Gid15, Gid16, Gid17, Gid18, Gid19,
    Gid20, Gid21, Gid22, Gid23, Gid24, Gid25, Gid26, Gid27, Gid28, Gid29,
    Gid30, Gid31, Gic0, Gic1, Gic2, Gic3, Gic4, Gic5, Gic6, Gic7, Gr;
  output God0, God1, God2, God3, God4, God5, God6, God7, God8, God9, God10,
    God11, God12, God13, God14, God15, God16, God17, God18, God19, God20,
    God21, God22, God23, God24, God25, God26, God27, God28, God29, God30,
    God31;
  wire n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n444, n445, n446, n447, n448, n450, n451,
    n452, n453, n454, n456, n457, n458, n459, n460, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n473, n474, n475, n476, n477, n479,
    n480, n481, n482, n483, n485, n486, n487, n488, n489, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n500, n501, n502, n504, n505, n506,
    n507, n508, n510, n511, n512, n513, n514, n516, n517, n518, n519, n520,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n532, n533, n534,
    n535, n536, n538, n539, n540, n541, n542, n544, n545, n546, n547, n548,
    n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568, n569, n571, n572, n573, n574,
    n575, n577, n578, n579, n580, n581, n583, n584, n585, n586, n587, n589,
    n590, n591, n592, n593, n594, n595, n596, n597, n598, n600, n601, n602,
    n603, n604, n606, n607, n608, n609, n610, n612, n613, n614, n615, n616,
    n618, n619, n620, n621, n622, n623, n624, n625, n627, n628, n629, n630,
    n631, n633, n634, n635, n636, n637, n639, n640, n641, n642, n643, n645,
    n646, n647, n648, n649, n650, n651, n653, n654, n655, n656, n657, n659,
    n660, n661, n662, n663, n665, n666, n667, n668, n669;
  inv1   g000(.a(Gic0), .O(n74));
  inv1   g001(.a(Gr), .O(n75));
  nor2   g002(.a(n75), .b(n74), .O(n76));
  inv1   g003(.a(n76), .O(n77));
  inv1   g004(.a(Gid16), .O(n78));
  nor2   g005(.a(Gid19), .b(n78), .O(n79));
  inv1   g006(.a(Gid19), .O(n80));
  nor2   g007(.a(n80), .b(Gid16), .O(n81));
  nor2   g008(.a(n81), .b(n79), .O(n82));
  inv1   g009(.a(n82), .O(n83));
  inv1   g010(.a(Gid17), .O(n84));
  nor2   g011(.a(Gid18), .b(n84), .O(n85));
  inv1   g012(.a(Gid18), .O(n86));
  nor2   g013(.a(n86), .b(Gid17), .O(n87));
  nor2   g014(.a(n87), .b(n85), .O(n88));
  nor2   g015(.a(n88), .b(n83), .O(n89));
  inv1   g016(.a(n88), .O(n90));
  nor2   g017(.a(n90), .b(n82), .O(n91));
  nor2   g018(.a(n91), .b(n89), .O(n92));
  inv1   g019(.a(n92), .O(n93));
  nor2   g020(.a(n93), .b(n77), .O(n94));
  nor2   g021(.a(n92), .b(n76), .O(n95));
  nor2   g022(.a(n95), .b(n94), .O(n96));
  inv1   g023(.a(n96), .O(n97));
  inv1   g024(.a(Gid0), .O(n98));
  nor2   g025(.a(Gid12), .b(n98), .O(n99));
  inv1   g026(.a(Gid12), .O(n100));
  nor2   g027(.a(n100), .b(Gid0), .O(n101));
  nor2   g028(.a(n101), .b(n99), .O(n102));
  inv1   g029(.a(n102), .O(n103));
  inv1   g030(.a(Gid4), .O(n104));
  nor2   g031(.a(Gid8), .b(n104), .O(n105));
  inv1   g032(.a(Gid8), .O(n106));
  nor2   g033(.a(n106), .b(Gid4), .O(n107));
  nor2   g034(.a(n107), .b(n105), .O(n108));
  nor2   g035(.a(n108), .b(n103), .O(n109));
  inv1   g036(.a(n108), .O(n110));
  nor2   g037(.a(n110), .b(n102), .O(n111));
  nor2   g038(.a(n111), .b(n109), .O(n112));
  inv1   g039(.a(n112), .O(n113));
  inv1   g040(.a(Gid20), .O(n114));
  nor2   g041(.a(Gid23), .b(n114), .O(n115));
  inv1   g042(.a(Gid23), .O(n116));
  nor2   g043(.a(n116), .b(Gid20), .O(n117));
  nor2   g044(.a(n117), .b(n115), .O(n118));
  inv1   g045(.a(n118), .O(n119));
  inv1   g046(.a(Gid21), .O(n120));
  nor2   g047(.a(Gid22), .b(n120), .O(n121));
  inv1   g048(.a(Gid22), .O(n122));
  nor2   g049(.a(n122), .b(Gid21), .O(n123));
  nor2   g050(.a(n123), .b(n121), .O(n124));
  nor2   g051(.a(n124), .b(n119), .O(n125));
  inv1   g052(.a(n124), .O(n126));
  nor2   g053(.a(n126), .b(n118), .O(n127));
  nor2   g054(.a(n127), .b(n125), .O(n128));
  nor2   g055(.a(n128), .b(n113), .O(n129));
  inv1   g056(.a(n128), .O(n130));
  nor2   g057(.a(n130), .b(n112), .O(n131));
  nor2   g058(.a(n131), .b(n129), .O(n132));
  inv1   g059(.a(n132), .O(n133));
  nor2   g060(.a(n133), .b(n97), .O(n134));
  nor2   g061(.a(n132), .b(n96), .O(n135));
  nor2   g062(.a(n135), .b(n134), .O(n136));
  inv1   g063(.a(n136), .O(n137));
  inv1   g064(.a(Gic7), .O(n138));
  nor2   g065(.a(n75), .b(n138), .O(n139));
  inv1   g066(.a(n139), .O(n140));
  nor2   g067(.a(Gid7), .b(n104), .O(n141));
  inv1   g068(.a(Gid7), .O(n142));
  nor2   g069(.a(n142), .b(Gid4), .O(n143));
  nor2   g070(.a(n143), .b(n141), .O(n144));
  inv1   g071(.a(n144), .O(n145));
  inv1   g072(.a(Gid5), .O(n146));
  nor2   g073(.a(Gid6), .b(n146), .O(n147));
  inv1   g074(.a(Gid6), .O(n148));
  nor2   g075(.a(n148), .b(Gid5), .O(n149));
  nor2   g076(.a(n149), .b(n147), .O(n150));
  nor2   g077(.a(n150), .b(n145), .O(n151));
  inv1   g078(.a(n150), .O(n152));
  nor2   g079(.a(n152), .b(n144), .O(n153));
  nor2   g080(.a(n153), .b(n151), .O(n154));
  inv1   g081(.a(n154), .O(n155));
  nor2   g082(.a(n155), .b(n140), .O(n156));
  nor2   g083(.a(n154), .b(n139), .O(n157));
  nor2   g084(.a(n157), .b(n156), .O(n158));
  inv1   g085(.a(n158), .O(n159));
  nor2   g086(.a(Gid15), .b(n100), .O(n160));
  inv1   g087(.a(Gid15), .O(n161));
  nor2   g088(.a(n161), .b(Gid12), .O(n162));
  nor2   g089(.a(n162), .b(n160), .O(n163));
  inv1   g090(.a(n163), .O(n164));
  inv1   g091(.a(Gid13), .O(n165));
  nor2   g092(.a(Gid14), .b(n165), .O(n166));
  inv1   g093(.a(Gid14), .O(n167));
  nor2   g094(.a(n167), .b(Gid13), .O(n168));
  nor2   g095(.a(n168), .b(n166), .O(n169));
  nor2   g096(.a(n169), .b(n164), .O(n170));
  inv1   g097(.a(n169), .O(n171));
  nor2   g098(.a(n171), .b(n163), .O(n172));
  nor2   g099(.a(n172), .b(n170), .O(n173));
  inv1   g100(.a(n173), .O(n174));
  nor2   g101(.a(Gid31), .b(n80), .O(n175));
  inv1   g102(.a(Gid31), .O(n176));
  nor2   g103(.a(n176), .b(Gid19), .O(n177));
  nor2   g104(.a(n177), .b(n175), .O(n178));
  inv1   g105(.a(n178), .O(n179));
  nor2   g106(.a(Gid27), .b(n116), .O(n180));
  inv1   g107(.a(Gid27), .O(n181));
  nor2   g108(.a(n181), .b(Gid23), .O(n182));
  nor2   g109(.a(n182), .b(n180), .O(n183));
  nor2   g110(.a(n183), .b(n179), .O(n184));
  inv1   g111(.a(n183), .O(n185));
  nor2   g112(.a(n185), .b(n178), .O(n186));
  nor2   g113(.a(n186), .b(n184), .O(n187));
  nor2   g114(.a(n187), .b(n174), .O(n188));
  inv1   g115(.a(n187), .O(n189));
  nor2   g116(.a(n189), .b(n173), .O(n190));
  nor2   g117(.a(n190), .b(n188), .O(n191));
  inv1   g118(.a(n191), .O(n192));
  nor2   g119(.a(n192), .b(n159), .O(n193));
  nor2   g120(.a(n191), .b(n158), .O(n194));
  nor2   g121(.a(n194), .b(n193), .O(n195));
  inv1   g122(.a(Gic6), .O(n196));
  nor2   g123(.a(n75), .b(n196), .O(n197));
  inv1   g124(.a(n197), .O(n198));
  nor2   g125(.a(Gid3), .b(n98), .O(n199));
  inv1   g126(.a(Gid3), .O(n200));
  nor2   g127(.a(n200), .b(Gid0), .O(n201));
  nor2   g128(.a(n201), .b(n199), .O(n202));
  inv1   g129(.a(n202), .O(n203));
  inv1   g130(.a(Gid1), .O(n204));
  nor2   g131(.a(Gid2), .b(n204), .O(n205));
  inv1   g132(.a(Gid2), .O(n206));
  nor2   g133(.a(n206), .b(Gid1), .O(n207));
  nor2   g134(.a(n207), .b(n205), .O(n208));
  nor2   g135(.a(n208), .b(n203), .O(n209));
  inv1   g136(.a(n208), .O(n210));
  nor2   g137(.a(n210), .b(n202), .O(n211));
  nor2   g138(.a(n211), .b(n209), .O(n212));
  inv1   g139(.a(n212), .O(n213));
  nor2   g140(.a(n213), .b(n198), .O(n214));
  nor2   g141(.a(n212), .b(n197), .O(n215));
  nor2   g142(.a(n215), .b(n214), .O(n216));
  inv1   g143(.a(n216), .O(n217));
  nor2   g144(.a(Gid11), .b(n106), .O(n218));
  inv1   g145(.a(Gid11), .O(n219));
  nor2   g146(.a(n219), .b(Gid8), .O(n220));
  nor2   g147(.a(n220), .b(n218), .O(n221));
  inv1   g148(.a(n221), .O(n222));
  inv1   g149(.a(Gid9), .O(n223));
  nor2   g150(.a(Gid10), .b(n223), .O(n224));
  inv1   g151(.a(Gid10), .O(n225));
  nor2   g152(.a(n225), .b(Gid9), .O(n226));
  nor2   g153(.a(n226), .b(n224), .O(n227));
  nor2   g154(.a(n227), .b(n222), .O(n228));
  inv1   g155(.a(n227), .O(n229));
  nor2   g156(.a(n229), .b(n221), .O(n230));
  nor2   g157(.a(n230), .b(n228), .O(n231));
  inv1   g158(.a(n231), .O(n232));
  nor2   g159(.a(Gid30), .b(n86), .O(n233));
  inv1   g160(.a(Gid30), .O(n234));
  nor2   g161(.a(n234), .b(Gid18), .O(n235));
  nor2   g162(.a(n235), .b(n233), .O(n236));
  inv1   g163(.a(n236), .O(n237));
  nor2   g164(.a(Gid26), .b(n122), .O(n238));
  inv1   g165(.a(Gid26), .O(n239));
  nor2   g166(.a(n239), .b(Gid22), .O(n240));
  nor2   g167(.a(n240), .b(n238), .O(n241));
  nor2   g168(.a(n241), .b(n237), .O(n242));
  inv1   g169(.a(n241), .O(n243));
  nor2   g170(.a(n243), .b(n236), .O(n244));
  nor2   g171(.a(n244), .b(n242), .O(n245));
  nor2   g172(.a(n245), .b(n232), .O(n246));
  inv1   g173(.a(n245), .O(n247));
  nor2   g174(.a(n247), .b(n231), .O(n248));
  nor2   g175(.a(n248), .b(n246), .O(n249));
  inv1   g176(.a(n249), .O(n250));
  nor2   g177(.a(n250), .b(n217), .O(n251));
  nor2   g178(.a(n249), .b(n216), .O(n252));
  nor2   g179(.a(n252), .b(n251), .O(n253));
  inv1   g180(.a(n253), .O(n254));
  nor2   g181(.a(n254), .b(n195), .O(n255));
  inv1   g182(.a(n255), .O(n256));
  inv1   g183(.a(Gic4), .O(n257));
  nor2   g184(.a(n75), .b(n257), .O(n258));
  inv1   g185(.a(n258), .O(n259));
  nor2   g186(.a(n259), .b(n155), .O(n260));
  nor2   g187(.a(n258), .b(n154), .O(n261));
  nor2   g188(.a(n261), .b(n260), .O(n262));
  inv1   g189(.a(n262), .O(n263));
  nor2   g190(.a(Gid28), .b(n78), .O(n264));
  inv1   g191(.a(Gid28), .O(n265));
  nor2   g192(.a(n265), .b(Gid16), .O(n266));
  nor2   g193(.a(n266), .b(n264), .O(n267));
  inv1   g194(.a(n267), .O(n268));
  nor2   g195(.a(Gid24), .b(n114), .O(n269));
  inv1   g196(.a(Gid24), .O(n270));
  nor2   g197(.a(n270), .b(Gid20), .O(n271));
  nor2   g198(.a(n271), .b(n269), .O(n272));
  nor2   g199(.a(n272), .b(n268), .O(n273));
  inv1   g200(.a(n272), .O(n274));
  nor2   g201(.a(n274), .b(n267), .O(n275));
  nor2   g202(.a(n275), .b(n273), .O(n276));
  nor2   g203(.a(n276), .b(n213), .O(n277));
  inv1   g204(.a(n276), .O(n278));
  nor2   g205(.a(n278), .b(n212), .O(n279));
  nor2   g206(.a(n279), .b(n277), .O(n280));
  inv1   g207(.a(n280), .O(n281));
  nor2   g208(.a(n281), .b(n263), .O(n282));
  nor2   g209(.a(n280), .b(n262), .O(n283));
  nor2   g210(.a(n283), .b(n282), .O(n284));
  inv1   g211(.a(n284), .O(n285));
  inv1   g212(.a(Gic5), .O(n286));
  nor2   g213(.a(n75), .b(n286), .O(n287));
  inv1   g214(.a(n287), .O(n288));
  nor2   g215(.a(n288), .b(n174), .O(n289));
  nor2   g216(.a(n287), .b(n173), .O(n290));
  nor2   g217(.a(n290), .b(n289), .O(n291));
  inv1   g218(.a(n291), .O(n292));
  nor2   g219(.a(Gid29), .b(n84), .O(n293));
  inv1   g220(.a(Gid29), .O(n294));
  nor2   g221(.a(n294), .b(Gid17), .O(n295));
  nor2   g222(.a(n295), .b(n293), .O(n296));
  inv1   g223(.a(n296), .O(n297));
  nor2   g224(.a(Gid25), .b(n120), .O(n298));
  inv1   g225(.a(Gid25), .O(n299));
  nor2   g226(.a(n299), .b(Gid21), .O(n300));
  nor2   g227(.a(n300), .b(n298), .O(n301));
  nor2   g228(.a(n301), .b(n297), .O(n302));
  inv1   g229(.a(n301), .O(n303));
  nor2   g230(.a(n303), .b(n296), .O(n304));
  nor2   g231(.a(n304), .b(n302), .O(n305));
  nor2   g232(.a(n305), .b(n232), .O(n306));
  inv1   g233(.a(n305), .O(n307));
  nor2   g234(.a(n307), .b(n231), .O(n308));
  nor2   g235(.a(n308), .b(n306), .O(n309));
  inv1   g236(.a(n309), .O(n310));
  nor2   g237(.a(n310), .b(n292), .O(n311));
  nor2   g238(.a(n309), .b(n291), .O(n312));
  nor2   g239(.a(n312), .b(n311), .O(n313));
  nor2   g240(.a(n313), .b(n285), .O(n314));
  inv1   g241(.a(n314), .O(n315));
  inv1   g242(.a(Gic1), .O(n316));
  nor2   g243(.a(n75), .b(n316), .O(n317));
  inv1   g244(.a(n317), .O(n318));
  nor2   g245(.a(Gid31), .b(n265), .O(n319));
  nor2   g246(.a(n176), .b(Gid28), .O(n320));
  nor2   g247(.a(n320), .b(n319), .O(n321));
  inv1   g248(.a(n321), .O(n322));
  nor2   g249(.a(Gid30), .b(n294), .O(n323));
  nor2   g250(.a(n234), .b(Gid29), .O(n324));
  nor2   g251(.a(n324), .b(n323), .O(n325));
  nor2   g252(.a(n325), .b(n322), .O(n326));
  inv1   g253(.a(n325), .O(n327));
  nor2   g254(.a(n327), .b(n321), .O(n328));
  nor2   g255(.a(n328), .b(n326), .O(n329));
  inv1   g256(.a(n329), .O(n330));
  nor2   g257(.a(n330), .b(n318), .O(n331));
  nor2   g258(.a(n329), .b(n317), .O(n332));
  nor2   g259(.a(n332), .b(n331), .O(n333));
  inv1   g260(.a(n333), .O(n334));
  nor2   g261(.a(Gid13), .b(n204), .O(n335));
  nor2   g262(.a(n165), .b(Gid1), .O(n336));
  nor2   g263(.a(n336), .b(n335), .O(n337));
  inv1   g264(.a(n337), .O(n338));
  nor2   g265(.a(Gid9), .b(n146), .O(n339));
  nor2   g266(.a(n223), .b(Gid5), .O(n340));
  nor2   g267(.a(n340), .b(n339), .O(n341));
  nor2   g268(.a(n341), .b(n338), .O(n342));
  inv1   g269(.a(n341), .O(n343));
  nor2   g270(.a(n343), .b(n337), .O(n344));
  nor2   g271(.a(n344), .b(n342), .O(n345));
  inv1   g272(.a(n345), .O(n346));
  nor2   g273(.a(Gid27), .b(n270), .O(n347));
  nor2   g274(.a(n181), .b(Gid24), .O(n348));
  nor2   g275(.a(n348), .b(n347), .O(n349));
  inv1   g276(.a(n349), .O(n350));
  nor2   g277(.a(Gid26), .b(n299), .O(n351));
  nor2   g278(.a(n239), .b(Gid25), .O(n352));
  nor2   g279(.a(n352), .b(n351), .O(n353));
  nor2   g280(.a(n353), .b(n350), .O(n354));
  inv1   g281(.a(n353), .O(n355));
  nor2   g282(.a(n355), .b(n349), .O(n356));
  nor2   g283(.a(n356), .b(n354), .O(n357));
  nor2   g284(.a(n357), .b(n346), .O(n358));
  inv1   g285(.a(n357), .O(n359));
  nor2   g286(.a(n359), .b(n345), .O(n360));
  nor2   g287(.a(n360), .b(n358), .O(n361));
  inv1   g288(.a(n361), .O(n362));
  nor2   g289(.a(n362), .b(n334), .O(n363));
  nor2   g290(.a(n361), .b(n333), .O(n364));
  nor2   g291(.a(n364), .b(n363), .O(n365));
  inv1   g292(.a(n365), .O(n366));
  nor2   g293(.a(n366), .b(n136), .O(n367));
  nor2   g294(.a(n365), .b(n137), .O(n368));
  nor2   g295(.a(n368), .b(n367), .O(n369));
  inv1   g296(.a(Gic2), .O(n370));
  nor2   g297(.a(n75), .b(n370), .O(n371));
  inv1   g298(.a(n371), .O(n372));
  nor2   g299(.a(n372), .b(n93), .O(n373));
  nor2   g300(.a(n371), .b(n92), .O(n374));
  nor2   g301(.a(n374), .b(n373), .O(n375));
  inv1   g302(.a(n375), .O(n376));
  nor2   g303(.a(Gid14), .b(n206), .O(n377));
  nor2   g304(.a(n167), .b(Gid2), .O(n378));
  nor2   g305(.a(n378), .b(n377), .O(n379));
  inv1   g306(.a(n379), .O(n380));
  nor2   g307(.a(Gid10), .b(n148), .O(n381));
  nor2   g308(.a(n225), .b(Gid6), .O(n382));
  nor2   g309(.a(n382), .b(n381), .O(n383));
  nor2   g310(.a(n383), .b(n380), .O(n384));
  inv1   g311(.a(n383), .O(n385));
  nor2   g312(.a(n385), .b(n379), .O(n386));
  nor2   g313(.a(n386), .b(n384), .O(n387));
  nor2   g314(.a(n387), .b(n359), .O(n388));
  inv1   g315(.a(n387), .O(n389));
  nor2   g316(.a(n389), .b(n357), .O(n390));
  nor2   g317(.a(n390), .b(n388), .O(n391));
  inv1   g318(.a(n391), .O(n392));
  nor2   g319(.a(n392), .b(n376), .O(n393));
  nor2   g320(.a(n391), .b(n375), .O(n394));
  nor2   g321(.a(n394), .b(n393), .O(n395));
  inv1   g322(.a(Gic3), .O(n396));
  nor2   g323(.a(n75), .b(n396), .O(n397));
  inv1   g324(.a(n397), .O(n398));
  nor2   g325(.a(n398), .b(n130), .O(n399));
  nor2   g326(.a(n397), .b(n128), .O(n400));
  nor2   g327(.a(n400), .b(n399), .O(n401));
  inv1   g328(.a(n401), .O(n402));
  nor2   g329(.a(Gid15), .b(n200), .O(n403));
  nor2   g330(.a(n161), .b(Gid3), .O(n404));
  nor2   g331(.a(n404), .b(n403), .O(n405));
  inv1   g332(.a(n405), .O(n406));
  nor2   g333(.a(Gid11), .b(n142), .O(n407));
  nor2   g334(.a(n219), .b(Gid7), .O(n408));
  nor2   g335(.a(n408), .b(n407), .O(n409));
  nor2   g336(.a(n409), .b(n406), .O(n410));
  inv1   g337(.a(n409), .O(n411));
  nor2   g338(.a(n411), .b(n405), .O(n412));
  nor2   g339(.a(n412), .b(n410), .O(n413));
  nor2   g340(.a(n413), .b(n330), .O(n414));
  inv1   g341(.a(n413), .O(n415));
  nor2   g342(.a(n415), .b(n329), .O(n416));
  nor2   g343(.a(n416), .b(n414), .O(n417));
  inv1   g344(.a(n417), .O(n418));
  nor2   g345(.a(n418), .b(n402), .O(n419));
  nor2   g346(.a(n417), .b(n401), .O(n420));
  nor2   g347(.a(n420), .b(n419), .O(n421));
  nor2   g348(.a(n421), .b(n395), .O(n422));
  inv1   g349(.a(n422), .O(n423));
  nor2   g350(.a(n423), .b(n369), .O(n424));
  inv1   g351(.a(n421), .O(n425));
  nor2   g352(.a(n425), .b(n395), .O(n426));
  inv1   g353(.a(n395), .O(n427));
  nor2   g354(.a(n421), .b(n427), .O(n428));
  nor2   g355(.a(n428), .b(n426), .O(n429));
  nor2   g356(.a(n365), .b(n136), .O(n430));
  inv1   g357(.a(n430), .O(n431));
  nor2   g358(.a(n431), .b(n429), .O(n432));
  nor2   g359(.a(n432), .b(n424), .O(n433));
  nor2   g360(.a(n433), .b(n315), .O(n434));
  inv1   g361(.a(n434), .O(n435));
  nor2   g362(.a(n435), .b(n256), .O(n436));
  inv1   g363(.a(n436), .O(n437));
  nor2   g364(.a(n437), .b(n137), .O(n438));
  inv1   g365(.a(n438), .O(n439));
  nor2   g366(.a(n439), .b(Gid0), .O(n440));
  nor2   g367(.a(n438), .b(n98), .O(n441));
  nor2   g368(.a(n441), .b(n440), .O(n442));
  inv1   g369(.a(n442), .O(God0));
  nor2   g370(.a(n437), .b(n366), .O(n444));
  inv1   g371(.a(n444), .O(n445));
  nor2   g372(.a(n445), .b(Gid1), .O(n446));
  nor2   g373(.a(n444), .b(n204), .O(n447));
  nor2   g374(.a(n447), .b(n446), .O(n448));
  inv1   g375(.a(n448), .O(God1));
  nor2   g376(.a(n437), .b(n427), .O(n450));
  inv1   g377(.a(n450), .O(n451));
  nor2   g378(.a(n451), .b(Gid2), .O(n452));
  nor2   g379(.a(n450), .b(n206), .O(n453));
  nor2   g380(.a(n453), .b(n452), .O(n454));
  inv1   g381(.a(n454), .O(God2));
  nor2   g382(.a(n437), .b(n425), .O(n456));
  inv1   g383(.a(n456), .O(n457));
  nor2   g384(.a(n457), .b(Gid3), .O(n458));
  nor2   g385(.a(n456), .b(n200), .O(n459));
  nor2   g386(.a(n459), .b(n458), .O(n460));
  inv1   g387(.a(n460), .O(God3));
  inv1   g388(.a(n195), .O(n462));
  nor2   g389(.a(n253), .b(n462), .O(n463));
  inv1   g390(.a(n463), .O(n464));
  nor2   g391(.a(n464), .b(n435), .O(n465));
  inv1   g392(.a(n465), .O(n466));
  nor2   g393(.a(n466), .b(n137), .O(n467));
  inv1   g394(.a(n467), .O(n468));
  nor2   g395(.a(n468), .b(Gid4), .O(n469));
  nor2   g396(.a(n467), .b(n104), .O(n470));
  nor2   g397(.a(n470), .b(n469), .O(n471));
  inv1   g398(.a(n471), .O(God4));
  nor2   g399(.a(n466), .b(n366), .O(n473));
  inv1   g400(.a(n473), .O(n474));
  nor2   g401(.a(n474), .b(Gid5), .O(n475));
  nor2   g402(.a(n473), .b(n146), .O(n476));
  nor2   g403(.a(n476), .b(n475), .O(n477));
  inv1   g404(.a(n477), .O(God5));
  nor2   g405(.a(n466), .b(n427), .O(n479));
  inv1   g406(.a(n479), .O(n480));
  nor2   g407(.a(n480), .b(Gid6), .O(n481));
  nor2   g408(.a(n479), .b(n148), .O(n482));
  nor2   g409(.a(n482), .b(n481), .O(n483));
  inv1   g410(.a(n483), .O(God6));
  nor2   g411(.a(n466), .b(n425), .O(n485));
  inv1   g412(.a(n485), .O(n486));
  nor2   g413(.a(n486), .b(Gid7), .O(n487));
  nor2   g414(.a(n485), .b(n142), .O(n488));
  nor2   g415(.a(n488), .b(n487), .O(n489));
  inv1   g416(.a(n489), .O(God7));
  inv1   g417(.a(n313), .O(n491));
  nor2   g418(.a(n491), .b(n284), .O(n492));
  inv1   g419(.a(n492), .O(n493));
  nor2   g420(.a(n493), .b(n256), .O(n494));
  inv1   g421(.a(n494), .O(n495));
  nor2   g422(.a(n495), .b(n433), .O(n496));
  inv1   g423(.a(n496), .O(n497));
  nor2   g424(.a(n497), .b(n137), .O(n498));
  inv1   g425(.a(n498), .O(n499));
  nor2   g426(.a(n499), .b(Gid8), .O(n500));
  nor2   g427(.a(n498), .b(n106), .O(n501));
  nor2   g428(.a(n501), .b(n500), .O(n502));
  inv1   g429(.a(n502), .O(God8));
  nor2   g430(.a(n497), .b(n366), .O(n504));
  inv1   g431(.a(n504), .O(n505));
  nor2   g432(.a(n505), .b(Gid9), .O(n506));
  nor2   g433(.a(n504), .b(n223), .O(n507));
  nor2   g434(.a(n507), .b(n506), .O(n508));
  inv1   g435(.a(n508), .O(God9));
  nor2   g436(.a(n497), .b(n427), .O(n510));
  inv1   g437(.a(n510), .O(n511));
  nor2   g438(.a(n511), .b(Gid10), .O(n512));
  nor2   g439(.a(n510), .b(n225), .O(n513));
  nor2   g440(.a(n513), .b(n512), .O(n514));
  inv1   g441(.a(n514), .O(God10));
  nor2   g442(.a(n497), .b(n425), .O(n516));
  inv1   g443(.a(n516), .O(n517));
  nor2   g444(.a(n517), .b(Gid11), .O(n518));
  nor2   g445(.a(n516), .b(n219), .O(n519));
  nor2   g446(.a(n519), .b(n518), .O(n520));
  inv1   g447(.a(n520), .O(God11));
  nor2   g448(.a(n493), .b(n464), .O(n522));
  inv1   g449(.a(n522), .O(n523));
  nor2   g450(.a(n523), .b(n433), .O(n524));
  inv1   g451(.a(n524), .O(n525));
  nor2   g452(.a(n525), .b(n137), .O(n526));
  inv1   g453(.a(n526), .O(n527));
  nor2   g454(.a(n527), .b(Gid12), .O(n528));
  nor2   g455(.a(n526), .b(n100), .O(n529));
  nor2   g456(.a(n529), .b(n528), .O(n530));
  inv1   g457(.a(n530), .O(God12));
  nor2   g458(.a(n525), .b(n366), .O(n532));
  inv1   g459(.a(n532), .O(n533));
  nor2   g460(.a(n533), .b(Gid13), .O(n534));
  nor2   g461(.a(n532), .b(n165), .O(n535));
  nor2   g462(.a(n535), .b(n534), .O(n536));
  inv1   g463(.a(n536), .O(God13));
  nor2   g464(.a(n525), .b(n427), .O(n538));
  inv1   g465(.a(n538), .O(n539));
  nor2   g466(.a(n539), .b(Gid14), .O(n540));
  nor2   g467(.a(n538), .b(n167), .O(n541));
  nor2   g468(.a(n541), .b(n540), .O(n542));
  inv1   g469(.a(n542), .O(God14));
  nor2   g470(.a(n525), .b(n425), .O(n544));
  inv1   g471(.a(n544), .O(n545));
  nor2   g472(.a(n545), .b(Gid15), .O(n546));
  nor2   g473(.a(n544), .b(n161), .O(n547));
  nor2   g474(.a(n547), .b(n546), .O(n548));
  inv1   g475(.a(n548), .O(God15));
  inv1   g476(.a(n368), .O(n550));
  inv1   g477(.a(n428), .O(n551));
  nor2   g478(.a(n463), .b(n255), .O(n552));
  nor2   g479(.a(n313), .b(n284), .O(n553));
  inv1   g480(.a(n553), .O(n554));
  nor2   g481(.a(n554), .b(n552), .O(n555));
  nor2   g482(.a(n492), .b(n314), .O(n556));
  nor2   g483(.a(n253), .b(n195), .O(n557));
  inv1   g484(.a(n557), .O(n558));
  nor2   g485(.a(n558), .b(n556), .O(n559));
  nor2   g486(.a(n559), .b(n555), .O(n560));
  nor2   g487(.a(n560), .b(n551), .O(n561));
  inv1   g488(.a(n561), .O(n562));
  nor2   g489(.a(n562), .b(n550), .O(n563));
  inv1   g490(.a(n563), .O(n564));
  nor2   g491(.a(n564), .b(n285), .O(n565));
  inv1   g492(.a(n565), .O(n566));
  nor2   g493(.a(n566), .b(Gid16), .O(n567));
  nor2   g494(.a(n565), .b(n78), .O(n568));
  nor2   g495(.a(n568), .b(n567), .O(n569));
  inv1   g496(.a(n569), .O(God16));
  nor2   g497(.a(n564), .b(n491), .O(n571));
  inv1   g498(.a(n571), .O(n572));
  nor2   g499(.a(n572), .b(Gid17), .O(n573));
  nor2   g500(.a(n571), .b(n84), .O(n574));
  nor2   g501(.a(n574), .b(n573), .O(n575));
  inv1   g502(.a(n575), .O(God17));
  nor2   g503(.a(n564), .b(n254), .O(n577));
  inv1   g504(.a(n577), .O(n578));
  nor2   g505(.a(n578), .b(Gid18), .O(n579));
  nor2   g506(.a(n577), .b(n86), .O(n580));
  nor2   g507(.a(n580), .b(n579), .O(n581));
  inv1   g508(.a(n581), .O(God18));
  nor2   g509(.a(n564), .b(n462), .O(n583));
  inv1   g510(.a(n583), .O(n584));
  nor2   g511(.a(n584), .b(Gid19), .O(n585));
  nor2   g512(.a(n583), .b(n80), .O(n586));
  nor2   g513(.a(n586), .b(n585), .O(n587));
  inv1   g514(.a(n587), .O(God19));
  inv1   g515(.a(n426), .O(n589));
  nor2   g516(.a(n560), .b(n589), .O(n590));
  inv1   g517(.a(n590), .O(n591));
  nor2   g518(.a(n591), .b(n550), .O(n592));
  inv1   g519(.a(n592), .O(n593));
  nor2   g520(.a(n593), .b(n285), .O(n594));
  inv1   g521(.a(n594), .O(n595));
  nor2   g522(.a(n595), .b(Gid20), .O(n596));
  nor2   g523(.a(n594), .b(n114), .O(n597));
  nor2   g524(.a(n597), .b(n596), .O(n598));
  inv1   g525(.a(n598), .O(God20));
  nor2   g526(.a(n593), .b(n491), .O(n600));
  inv1   g527(.a(n600), .O(n601));
  nor2   g528(.a(n601), .b(Gid21), .O(n602));
  nor2   g529(.a(n600), .b(n120), .O(n603));
  nor2   g530(.a(n603), .b(n602), .O(n604));
  inv1   g531(.a(n604), .O(God21));
  nor2   g532(.a(n593), .b(n254), .O(n606));
  inv1   g533(.a(n606), .O(n607));
  nor2   g534(.a(n607), .b(Gid22), .O(n608));
  nor2   g535(.a(n606), .b(n122), .O(n609));
  nor2   g536(.a(n609), .b(n608), .O(n610));
  inv1   g537(.a(n610), .O(God22));
  nor2   g538(.a(n593), .b(n462), .O(n612));
  inv1   g539(.a(n612), .O(n613));
  nor2   g540(.a(n613), .b(Gid23), .O(n614));
  nor2   g541(.a(n612), .b(n116), .O(n615));
  nor2   g542(.a(n615), .b(n614), .O(n616));
  inv1   g543(.a(n616), .O(God23));
  inv1   g544(.a(n367), .O(n618));
  nor2   g545(.a(n562), .b(n618), .O(n619));
  inv1   g546(.a(n619), .O(n620));
  nor2   g547(.a(n620), .b(n285), .O(n621));
  inv1   g548(.a(n621), .O(n622));
  nor2   g549(.a(n622), .b(Gid24), .O(n623));
  nor2   g550(.a(n621), .b(n270), .O(n624));
  nor2   g551(.a(n624), .b(n623), .O(n625));
  inv1   g552(.a(n625), .O(God24));
  nor2   g553(.a(n620), .b(n491), .O(n627));
  inv1   g554(.a(n627), .O(n628));
  nor2   g555(.a(n628), .b(Gid25), .O(n629));
  nor2   g556(.a(n627), .b(n299), .O(n630));
  nor2   g557(.a(n630), .b(n629), .O(n631));
  inv1   g558(.a(n631), .O(God25));
  nor2   g559(.a(n620), .b(n254), .O(n633));
  inv1   g560(.a(n633), .O(n634));
  nor2   g561(.a(n634), .b(Gid26), .O(n635));
  nor2   g562(.a(n633), .b(n239), .O(n636));
  nor2   g563(.a(n636), .b(n635), .O(n637));
  inv1   g564(.a(n637), .O(God26));
  nor2   g565(.a(n620), .b(n462), .O(n639));
  inv1   g566(.a(n639), .O(n640));
  nor2   g567(.a(n640), .b(Gid27), .O(n641));
  nor2   g568(.a(n639), .b(n181), .O(n642));
  nor2   g569(.a(n642), .b(n641), .O(n643));
  inv1   g570(.a(n643), .O(God27));
  nor2   g571(.a(n591), .b(n618), .O(n645));
  inv1   g572(.a(n645), .O(n646));
  nor2   g573(.a(n646), .b(n285), .O(n647));
  inv1   g574(.a(n647), .O(n648));
  nor2   g575(.a(n648), .b(Gid28), .O(n649));
  nor2   g576(.a(n647), .b(n265), .O(n650));
  nor2   g577(.a(n650), .b(n649), .O(n651));
  inv1   g578(.a(n651), .O(God28));
  nor2   g579(.a(n646), .b(n491), .O(n653));
  inv1   g580(.a(n653), .O(n654));
  nor2   g581(.a(n654), .b(Gid29), .O(n655));
  nor2   g582(.a(n653), .b(n294), .O(n656));
  nor2   g583(.a(n656), .b(n655), .O(n657));
  inv1   g584(.a(n657), .O(God29));
  nor2   g585(.a(n646), .b(n254), .O(n659));
  inv1   g586(.a(n659), .O(n660));
  nor2   g587(.a(n660), .b(Gid30), .O(n661));
  nor2   g588(.a(n659), .b(n234), .O(n662));
  nor2   g589(.a(n662), .b(n661), .O(n663));
  inv1   g590(.a(n663), .O(God30));
  nor2   g591(.a(n646), .b(n462), .O(n665));
  inv1   g592(.a(n665), .O(n666));
  nor2   g593(.a(n666), .b(Gid31), .O(n667));
  nor2   g594(.a(n665), .b(n176), .O(n668));
  nor2   g595(.a(n668), .b(n667), .O(n669));
  inv1   g596(.a(n669), .O(God31));
endmodule


