// Benchmark "c1908_blif" written by ABC on Sun Mar 24 18:39:13 2019

module c1908_blif  ( 
    G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
    G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237,
    G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n359, n360, n361, n362, n363, n364, n365, n366,
    n367, n369, n370, n371, n372, n373, n374, n375, n376, n377, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n395, n396, n397, n398, n399, n400, n401, n402, n403, n405, n406,
    n407, n408, n409, n410, n411, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n426, n427, n428, n429, n430, n432, n433,
    n434, n435, n436, n437, n438, n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n452, n453, n454, n455, n456, n457, n458, n460,
    n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n473,
    n474, n475, n476, n477, n479, n480, n481, n482, n483, n484, n485, n486,
    n487, n489, n490, n491, n492, n493, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n560, n561,
    n562, n563, n564, n565, n566, n567, n568, n570, n571, n572, n573, n574,
    n575, n576, n577, n579, n580, n581, n582, n583, n584, n585, n586, n588,
    n589, n590, n591, n592, n593, n594, n595, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n607, n608, n609, n610, n611, n612, n613, n614,
    n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
    n628, n630, n631, n632, n633, n634, n635, n636, n637;
  inv1   g000(.a(G101), .O(n59));
  inv1   g001(.a(G110), .O(n60));
  inv1   g002(.a(G137), .O(n61));
  inv1   g003(.a(G119), .O(n62));
  nor2   g004(.a(G128), .b(n62), .O(n63));
  inv1   g005(.a(G128), .O(n64));
  nor2   g006(.a(n64), .b(G119), .O(n65));
  nor2   g007(.a(n65), .b(n63), .O(n66));
  inv1   g008(.a(n66), .O(n67));
  nor2   g009(.a(n67), .b(n61), .O(n68));
  nor2   g010(.a(n66), .b(G137), .O(n69));
  nor2   g011(.a(n69), .b(n68), .O(n70));
  nor2   g012(.a(n70), .b(n60), .O(n71));
  inv1   g013(.a(n70), .O(n72));
  nor2   g014(.a(n72), .b(G110), .O(n73));
  nor2   g015(.a(n73), .b(n71), .O(n74));
  inv1   g016(.a(n74), .O(n75));
  inv1   g017(.a(G221), .O(n76));
  inv1   g018(.a(G234), .O(n77));
  nor2   g019(.a(n77), .b(n76), .O(n78));
  inv1   g020(.a(n78), .O(n79));
  nor2   g021(.a(n79), .b(G953), .O(n80));
  inv1   g022(.a(n80), .O(n81));
  inv1   g023(.a(G146), .O(n82));
  inv1   g024(.a(G125), .O(n83));
  nor2   g025(.a(G140), .b(n83), .O(n84));
  inv1   g026(.a(G140), .O(n85));
  nor2   g027(.a(n85), .b(G125), .O(n86));
  nor2   g028(.a(n86), .b(n84), .O(n87));
  nor2   g029(.a(n87), .b(n82), .O(n88));
  inv1   g030(.a(n87), .O(n89));
  nor2   g031(.a(n89), .b(G146), .O(n90));
  nor2   g032(.a(n90), .b(n88), .O(n91));
  nor2   g033(.a(n91), .b(n81), .O(n92));
  inv1   g034(.a(n91), .O(n93));
  nor2   g035(.a(n93), .b(n80), .O(n94));
  nor2   g036(.a(n94), .b(n92), .O(n95));
  inv1   g037(.a(n95), .O(n96));
  nor2   g038(.a(n96), .b(n75), .O(n97));
  nor2   g039(.a(n95), .b(n74), .O(n98));
  nor2   g040(.a(n98), .b(n97), .O(n99));
  nor2   g041(.a(n99), .b(G902), .O(n100));
  inv1   g042(.a(G217), .O(n101));
  nor2   g043(.a(G902), .b(n77), .O(n102));
  nor2   g044(.a(n102), .b(n101), .O(n103));
  inv1   g045(.a(n103), .O(n104));
  nor2   g046(.a(n104), .b(n100), .O(n105));
  inv1   g047(.a(n100), .O(n106));
  nor2   g048(.a(n103), .b(n106), .O(n107));
  nor2   g049(.a(n107), .b(n105), .O(n108));
  inv1   g050(.a(n108), .O(n109));
  inv1   g051(.a(G472), .O(n110));
  inv1   g052(.a(G113), .O(n111));
  inv1   g053(.a(G116), .O(n112));
  nor2   g054(.a(G119), .b(n112), .O(n113));
  nor2   g055(.a(n62), .b(G116), .O(n114));
  nor2   g056(.a(n114), .b(n113), .O(n115));
  nor2   g057(.a(n115), .b(n111), .O(n116));
  inv1   g058(.a(n115), .O(n117));
  nor2   g059(.a(n117), .b(G113), .O(n118));
  nor2   g060(.a(n118), .b(n116), .O(n119));
  inv1   g061(.a(n119), .O(n120));
  inv1   g062(.a(G210), .O(n121));
  nor2   g063(.a(G237), .b(n121), .O(n122));
  inv1   g064(.a(n122), .O(n123));
  nor2   g065(.a(n123), .b(G953), .O(n124));
  nor2   g066(.a(n124), .b(n59), .O(n125));
  inv1   g067(.a(n124), .O(n126));
  nor2   g068(.a(n126), .b(G101), .O(n127));
  nor2   g069(.a(n127), .b(n125), .O(n128));
  inv1   g070(.a(n128), .O(n129));
  inv1   g071(.a(G143), .O(n130));
  nor2   g072(.a(G146), .b(n130), .O(n131));
  nor2   g073(.a(n82), .b(G143), .O(n132));
  nor2   g074(.a(n132), .b(n131), .O(n133));
  nor2   g075(.a(n133), .b(n64), .O(n134));
  inv1   g076(.a(n133), .O(n135));
  nor2   g077(.a(n135), .b(G128), .O(n136));
  nor2   g078(.a(n136), .b(n134), .O(n137));
  inv1   g079(.a(n137), .O(n138));
  inv1   g080(.a(G131), .O(n139));
  inv1   g081(.a(G134), .O(n140));
  nor2   g082(.a(G137), .b(n140), .O(n141));
  nor2   g083(.a(n61), .b(G134), .O(n142));
  nor2   g084(.a(n142), .b(n141), .O(n143));
  nor2   g085(.a(n143), .b(n139), .O(n144));
  inv1   g086(.a(n143), .O(n145));
  nor2   g087(.a(n145), .b(G131), .O(n146));
  nor2   g088(.a(n146), .b(n144), .O(n147));
  inv1   g089(.a(n147), .O(n148));
  nor2   g090(.a(n148), .b(n138), .O(n149));
  nor2   g091(.a(n147), .b(n137), .O(n150));
  nor2   g092(.a(n150), .b(n149), .O(n151));
  nor2   g093(.a(n151), .b(n129), .O(n152));
  inv1   g094(.a(n151), .O(n153));
  nor2   g095(.a(n153), .b(n128), .O(n154));
  nor2   g096(.a(n154), .b(n152), .O(n155));
  inv1   g097(.a(n155), .O(n156));
  nor2   g098(.a(n156), .b(n120), .O(n157));
  nor2   g099(.a(n155), .b(n119), .O(n158));
  nor2   g100(.a(n158), .b(n157), .O(n159));
  inv1   g101(.a(n159), .O(n160));
  nor2   g102(.a(n160), .b(G902), .O(n161));
  nor2   g103(.a(n161), .b(n110), .O(n162));
  inv1   g104(.a(n161), .O(n163));
  nor2   g105(.a(n163), .b(G472), .O(n164));
  nor2   g106(.a(n164), .b(n162), .O(n165));
  nor2   g107(.a(n165), .b(n109), .O(n166));
  inv1   g108(.a(n166), .O(n167));
  inv1   g109(.a(G214), .O(n168));
  nor2   g110(.a(G902), .b(G237), .O(n169));
  nor2   g111(.a(n169), .b(n168), .O(n170));
  nor2   g112(.a(n169), .b(n121), .O(n171));
  nor2   g113(.a(G122), .b(n60), .O(n172));
  inv1   g114(.a(G122), .O(n173));
  nor2   g115(.a(n173), .b(G110), .O(n174));
  nor2   g116(.a(n174), .b(n172), .O(n175));
  inv1   g117(.a(n175), .O(n176));
  inv1   g118(.a(G104), .O(n177));
  nor2   g119(.a(G107), .b(n177), .O(n178));
  inv1   g120(.a(G107), .O(n179));
  nor2   g121(.a(n179), .b(G104), .O(n180));
  nor2   g122(.a(n180), .b(n178), .O(n181));
  nor2   g123(.a(n181), .b(n59), .O(n182));
  inv1   g124(.a(n181), .O(n183));
  nor2   g125(.a(n183), .b(G101), .O(n184));
  nor2   g126(.a(n184), .b(n182), .O(n185));
  nor2   g127(.a(n185), .b(n120), .O(n186));
  inv1   g128(.a(n185), .O(n187));
  nor2   g129(.a(n187), .b(n119), .O(n188));
  nor2   g130(.a(n188), .b(n186), .O(n189));
  inv1   g131(.a(n189), .O(n190));
  nor2   g132(.a(n190), .b(n176), .O(n191));
  nor2   g133(.a(n189), .b(n175), .O(n192));
  nor2   g134(.a(n192), .b(n191), .O(n193));
  inv1   g135(.a(n193), .O(n194));
  inv1   g136(.a(G224), .O(n195));
  nor2   g137(.a(G953), .b(n195), .O(n196));
  inv1   g138(.a(n196), .O(n197));
  nor2   g139(.a(n137), .b(n83), .O(n198));
  nor2   g140(.a(n138), .b(G125), .O(n199));
  nor2   g141(.a(n199), .b(n198), .O(n200));
  nor2   g142(.a(n200), .b(n197), .O(n201));
  inv1   g143(.a(n200), .O(n202));
  nor2   g144(.a(n202), .b(n196), .O(n203));
  nor2   g145(.a(n203), .b(n201), .O(n204));
  inv1   g146(.a(n204), .O(n205));
  nor2   g147(.a(n205), .b(n194), .O(n206));
  nor2   g148(.a(n204), .b(n193), .O(n207));
  nor2   g149(.a(n207), .b(n206), .O(n208));
  inv1   g150(.a(n208), .O(n209));
  nor2   g151(.a(n209), .b(G902), .O(n210));
  inv1   g152(.a(n210), .O(n211));
  nor2   g153(.a(n211), .b(n171), .O(n212));
  inv1   g154(.a(n171), .O(n213));
  nor2   g155(.a(n210), .b(n213), .O(n214));
  nor2   g156(.a(n214), .b(n212), .O(n215));
  nor2   g157(.a(n215), .b(n170), .O(n216));
  inv1   g158(.a(n216), .O(n217));
  nor2   g159(.a(n102), .b(n76), .O(n218));
  inv1   g160(.a(G469), .O(n219));
  inv1   g161(.a(G227), .O(n220));
  nor2   g162(.a(G953), .b(n220), .O(n221));
  nor2   g163(.a(n221), .b(n187), .O(n222));
  inv1   g164(.a(n221), .O(n223));
  nor2   g165(.a(n223), .b(n185), .O(n224));
  nor2   g166(.a(n224), .b(n222), .O(n225));
  inv1   g167(.a(n225), .O(n226));
  nor2   g168(.a(G140), .b(G110), .O(n227));
  nor2   g169(.a(n85), .b(n60), .O(n228));
  nor2   g170(.a(n228), .b(n227), .O(n229));
  inv1   g171(.a(n229), .O(n230));
  nor2   g172(.a(n230), .b(n151), .O(n231));
  nor2   g173(.a(n229), .b(n153), .O(n232));
  nor2   g174(.a(n232), .b(n231), .O(n233));
  inv1   g175(.a(n233), .O(n234));
  nor2   g176(.a(n234), .b(n226), .O(n235));
  nor2   g177(.a(n233), .b(n225), .O(n236));
  nor2   g178(.a(n236), .b(n235), .O(n237));
  inv1   g179(.a(n237), .O(n238));
  nor2   g180(.a(n238), .b(G902), .O(n239));
  nor2   g181(.a(n239), .b(n219), .O(n240));
  inv1   g182(.a(n239), .O(n241));
  nor2   g183(.a(n241), .b(G469), .O(n242));
  nor2   g184(.a(n242), .b(n240), .O(n243));
  nor2   g185(.a(n243), .b(n218), .O(n244));
  inv1   g186(.a(n244), .O(n245));
  nor2   g187(.a(n245), .b(n217), .O(n246));
  inv1   g188(.a(n246), .O(n247));
  nor2   g189(.a(n247), .b(n167), .O(n248));
  inv1   g190(.a(n248), .O(n249));
  inv1   g191(.a(G478), .O(n250));
  nor2   g192(.a(G134), .b(n179), .O(n251));
  nor2   g193(.a(n140), .b(G107), .O(n252));
  nor2   g194(.a(n252), .b(n251), .O(n253));
  inv1   g195(.a(n253), .O(n254));
  nor2   g196(.a(n77), .b(n101), .O(n255));
  inv1   g197(.a(n255), .O(n256));
  nor2   g198(.a(n256), .b(G953), .O(n257));
  nor2   g199(.a(n257), .b(n173), .O(n258));
  inv1   g200(.a(n257), .O(n259));
  nor2   g201(.a(n259), .b(G122), .O(n260));
  nor2   g202(.a(n260), .b(n258), .O(n261));
  inv1   g203(.a(n261), .O(n262));
  nor2   g204(.a(G143), .b(n64), .O(n263));
  nor2   g205(.a(n130), .b(G128), .O(n264));
  nor2   g206(.a(n264), .b(n263), .O(n265));
  inv1   g207(.a(n265), .O(n266));
  nor2   g208(.a(n266), .b(n112), .O(n267));
  nor2   g209(.a(n265), .b(G116), .O(n268));
  nor2   g210(.a(n268), .b(n267), .O(n269));
  nor2   g211(.a(n269), .b(n262), .O(n270));
  inv1   g212(.a(n269), .O(n271));
  nor2   g213(.a(n271), .b(n261), .O(n272));
  nor2   g214(.a(n272), .b(n270), .O(n273));
  inv1   g215(.a(n273), .O(n274));
  nor2   g216(.a(n274), .b(n254), .O(n275));
  nor2   g217(.a(n273), .b(n253), .O(n276));
  nor2   g218(.a(n276), .b(n275), .O(n277));
  inv1   g219(.a(n277), .O(n278));
  nor2   g220(.a(n278), .b(G902), .O(n279));
  nor2   g221(.a(n279), .b(n250), .O(n280));
  inv1   g222(.a(n279), .O(n281));
  nor2   g223(.a(n281), .b(G478), .O(n282));
  nor2   g224(.a(n282), .b(n280), .O(n283));
  inv1   g225(.a(n283), .O(n284));
  inv1   g226(.a(G475), .O(n285));
  nor2   g227(.a(G122), .b(n111), .O(n286));
  nor2   g228(.a(n173), .b(G113), .O(n287));
  nor2   g229(.a(n287), .b(n286), .O(n288));
  inv1   g230(.a(n288), .O(n289));
  nor2   g231(.a(n91), .b(n177), .O(n290));
  nor2   g232(.a(n93), .b(G104), .O(n291));
  nor2   g233(.a(n291), .b(n290), .O(n292));
  inv1   g234(.a(n292), .O(n293));
  nor2   g235(.a(n293), .b(n289), .O(n294));
  nor2   g236(.a(n292), .b(n288), .O(n295));
  nor2   g237(.a(n295), .b(n294), .O(n296));
  inv1   g238(.a(n296), .O(n297));
  nor2   g239(.a(G237), .b(n168), .O(n298));
  inv1   g240(.a(n298), .O(n299));
  nor2   g241(.a(n299), .b(G953), .O(n300));
  inv1   g242(.a(n300), .O(n301));
  nor2   g243(.a(G143), .b(n139), .O(n302));
  nor2   g244(.a(n130), .b(G131), .O(n303));
  nor2   g245(.a(n303), .b(n302), .O(n304));
  nor2   g246(.a(n304), .b(n301), .O(n305));
  inv1   g247(.a(n304), .O(n306));
  nor2   g248(.a(n306), .b(n300), .O(n307));
  nor2   g249(.a(n307), .b(n305), .O(n308));
  inv1   g250(.a(n308), .O(n309));
  nor2   g251(.a(n309), .b(n297), .O(n310));
  nor2   g252(.a(n308), .b(n296), .O(n311));
  nor2   g253(.a(n311), .b(n310), .O(n312));
  inv1   g254(.a(n312), .O(n313));
  nor2   g255(.a(n313), .b(G902), .O(n314));
  nor2   g256(.a(n314), .b(n285), .O(n315));
  inv1   g257(.a(n314), .O(n316));
  nor2   g258(.a(n316), .b(G475), .O(n317));
  nor2   g259(.a(n317), .b(n315), .O(n318));
  inv1   g260(.a(n318), .O(n319));
  nor2   g261(.a(n319), .b(n284), .O(n320));
  inv1   g262(.a(n320), .O(n321));
  inv1   g263(.a(G237), .O(n322));
  nor2   g264(.a(n322), .b(n77), .O(n323));
  inv1   g265(.a(G952), .O(n324));
  nor2   g266(.a(G953), .b(n324), .O(n325));
  inv1   g267(.a(n325), .O(n326));
  nor2   g268(.a(n326), .b(n323), .O(n327));
  inv1   g269(.a(G953), .O(n328));
  nor2   g270(.a(n328), .b(G898), .O(n329));
  inv1   g271(.a(n329), .O(n330));
  inv1   g272(.a(G902), .O(n331));
  nor2   g273(.a(n323), .b(n331), .O(n332));
  inv1   g274(.a(n332), .O(n333));
  nor2   g275(.a(n333), .b(n330), .O(n334));
  nor2   g276(.a(n334), .b(n327), .O(n335));
  nor2   g277(.a(n335), .b(n321), .O(n336));
  inv1   g278(.a(n336), .O(n337));
  nor2   g279(.a(n337), .b(n249), .O(n338));
  nor2   g280(.a(n338), .b(n59), .O(n339));
  inv1   g281(.a(n338), .O(n340));
  nor2   g282(.a(n340), .b(G101), .O(n341));
  nor2   g283(.a(n341), .b(n339), .O(n342));
  inv1   g284(.a(n342), .O(G3));
  inv1   g285(.a(n165), .O(n344));
  nor2   g286(.a(n344), .b(n109), .O(n345));
  inv1   g287(.a(n345), .O(n346));
  nor2   g288(.a(n346), .b(n247), .O(n347));
  inv1   g289(.a(n347), .O(n348));
  nor2   g290(.a(n318), .b(n284), .O(n349));
  inv1   g291(.a(n349), .O(n350));
  nor2   g292(.a(n350), .b(n335), .O(n351));
  inv1   g293(.a(n351), .O(n352));
  nor2   g294(.a(n352), .b(n348), .O(n353));
  nor2   g295(.a(n353), .b(n177), .O(n354));
  inv1   g296(.a(n353), .O(n355));
  nor2   g297(.a(n355), .b(G104), .O(n356));
  nor2   g298(.a(n356), .b(n354), .O(n357));
  inv1   g299(.a(n357), .O(G6));
  nor2   g300(.a(n319), .b(n283), .O(n359));
  inv1   g301(.a(n359), .O(n360));
  nor2   g302(.a(n360), .b(n335), .O(n361));
  inv1   g303(.a(n361), .O(n362));
  nor2   g304(.a(n362), .b(n348), .O(n363));
  nor2   g305(.a(n363), .b(n179), .O(n364));
  inv1   g306(.a(n363), .O(n365));
  nor2   g307(.a(n365), .b(G107), .O(n366));
  nor2   g308(.a(n366), .b(n364), .O(n367));
  inv1   g309(.a(n367), .O(G9));
  nor2   g310(.a(n344), .b(n108), .O(n369));
  inv1   g311(.a(n369), .O(n370));
  nor2   g312(.a(n370), .b(n247), .O(n371));
  inv1   g313(.a(n371), .O(n372));
  nor2   g314(.a(n372), .b(n337), .O(n373));
  nor2   g315(.a(n373), .b(n60), .O(n374));
  inv1   g316(.a(n373), .O(n375));
  nor2   g317(.a(n375), .b(G110), .O(n376));
  nor2   g318(.a(n376), .b(n374), .O(n377));
  inv1   g319(.a(n377), .O(G12));
  nor2   g320(.a(n165), .b(n108), .O(n379));
  inv1   g321(.a(n379), .O(n380));
  nor2   g322(.a(n380), .b(n247), .O(n381));
  inv1   g323(.a(n381), .O(n382));
  nor2   g324(.a(n328), .b(G900), .O(n383));
  inv1   g325(.a(n383), .O(n384));
  nor2   g326(.a(n384), .b(n333), .O(n385));
  nor2   g327(.a(n385), .b(n327), .O(n386));
  nor2   g328(.a(n386), .b(n360), .O(n387));
  inv1   g329(.a(n387), .O(n388));
  nor2   g330(.a(n388), .b(n382), .O(n389));
  nor2   g331(.a(n389), .b(n64), .O(n390));
  inv1   g332(.a(n389), .O(n391));
  nor2   g333(.a(n391), .b(G128), .O(n392));
  nor2   g334(.a(n392), .b(n390), .O(n393));
  inv1   g335(.a(n393), .O(G30));
  nor2   g336(.a(n318), .b(n283), .O(n395));
  inv1   g337(.a(n395), .O(n396));
  nor2   g338(.a(n396), .b(n386), .O(n397));
  inv1   g339(.a(n397), .O(n398));
  nor2   g340(.a(n398), .b(n249), .O(n399));
  nor2   g341(.a(n399), .b(n130), .O(n400));
  inv1   g342(.a(n399), .O(n401));
  nor2   g343(.a(n401), .b(G143), .O(n402));
  nor2   g344(.a(n402), .b(n400), .O(n403));
  inv1   g345(.a(n403), .O(G45));
  nor2   g346(.a(n386), .b(n350), .O(n405));
  inv1   g347(.a(n405), .O(n406));
  nor2   g348(.a(n406), .b(n382), .O(n407));
  nor2   g349(.a(n407), .b(n82), .O(n408));
  inv1   g350(.a(n407), .O(n409));
  nor2   g351(.a(n409), .b(G146), .O(n410));
  nor2   g352(.a(n410), .b(n408), .O(n411));
  inv1   g353(.a(n411), .O(G48));
  inv1   g354(.a(n243), .O(n413));
  nor2   g355(.a(n413), .b(n218), .O(n414));
  inv1   g356(.a(n414), .O(n415));
  nor2   g357(.a(n415), .b(n217), .O(n416));
  inv1   g358(.a(n416), .O(n417));
  nor2   g359(.a(n417), .b(n167), .O(n418));
  inv1   g360(.a(n418), .O(n419));
  nor2   g361(.a(n419), .b(n352), .O(n420));
  nor2   g362(.a(n420), .b(n111), .O(n421));
  inv1   g363(.a(n420), .O(n422));
  nor2   g364(.a(n422), .b(G113), .O(n423));
  nor2   g365(.a(n423), .b(n421), .O(n424));
  inv1   g366(.a(n424), .O(G15));
  nor2   g367(.a(n419), .b(n362), .O(n426));
  nor2   g368(.a(n426), .b(n112), .O(n427));
  inv1   g369(.a(n426), .O(n428));
  nor2   g370(.a(n428), .b(G116), .O(n429));
  nor2   g371(.a(n429), .b(n427), .O(n430));
  inv1   g372(.a(n430), .O(G18));
  nor2   g373(.a(n380), .b(n337), .O(n432));
  inv1   g374(.a(n432), .O(n433));
  nor2   g375(.a(n433), .b(n417), .O(n434));
  nor2   g376(.a(n434), .b(n62), .O(n435));
  inv1   g377(.a(n434), .O(n436));
  nor2   g378(.a(n436), .b(G119), .O(n437));
  nor2   g379(.a(n437), .b(n435), .O(n438));
  inv1   g380(.a(n438), .O(G21));
  nor2   g381(.a(n415), .b(n346), .O(n440));
  inv1   g382(.a(n440), .O(n441));
  nor2   g383(.a(n441), .b(n217), .O(n442));
  inv1   g384(.a(n442), .O(n443));
  nor2   g385(.a(n396), .b(n335), .O(n444));
  inv1   g386(.a(n444), .O(n445));
  nor2   g387(.a(n445), .b(n443), .O(n446));
  nor2   g388(.a(n446), .b(n173), .O(n447));
  inv1   g389(.a(n446), .O(n448));
  nor2   g390(.a(n448), .b(G122), .O(n449));
  nor2   g391(.a(n449), .b(n447), .O(n450));
  inv1   g392(.a(n450), .O(G24));
  nor2   g393(.a(n406), .b(n370), .O(n452));
  inv1   g394(.a(n452), .O(n453));
  nor2   g395(.a(n453), .b(n417), .O(n454));
  nor2   g396(.a(n454), .b(n83), .O(n455));
  inv1   g397(.a(n454), .O(n456));
  nor2   g398(.a(n456), .b(G125), .O(n457));
  nor2   g399(.a(n457), .b(n455), .O(n458));
  inv1   g400(.a(n458), .O(G27));
  inv1   g401(.a(n215), .O(n460));
  nor2   g402(.a(n460), .b(n170), .O(n461));
  inv1   g403(.a(n461), .O(n462));
  nor2   g404(.a(n462), .b(n245), .O(n463));
  inv1   g405(.a(n463), .O(n464));
  nor2   g406(.a(n464), .b(n167), .O(n465));
  inv1   g407(.a(n465), .O(n466));
  nor2   g408(.a(n466), .b(n406), .O(n467));
  nor2   g409(.a(n467), .b(n139), .O(n468));
  inv1   g410(.a(n467), .O(n469));
  nor2   g411(.a(n469), .b(G131), .O(n470));
  nor2   g412(.a(n470), .b(n468), .O(n471));
  inv1   g413(.a(n471), .O(G33));
  nor2   g414(.a(n466), .b(n388), .O(n473));
  nor2   g415(.a(n473), .b(n140), .O(n474));
  inv1   g416(.a(n473), .O(n475));
  nor2   g417(.a(n475), .b(G134), .O(n476));
  nor2   g418(.a(n476), .b(n474), .O(n477));
  inv1   g419(.a(n477), .O(G36));
  nor2   g420(.a(n386), .b(n321), .O(n479));
  inv1   g421(.a(n479), .O(n480));
  nor2   g422(.a(n480), .b(n380), .O(n481));
  inv1   g423(.a(n481), .O(n482));
  nor2   g424(.a(n482), .b(n464), .O(n483));
  nor2   g425(.a(n483), .b(n61), .O(n484));
  inv1   g426(.a(n483), .O(n485));
  nor2   g427(.a(n485), .b(G137), .O(n486));
  nor2   g428(.a(n486), .b(n484), .O(n487));
  inv1   g429(.a(n487), .O(G39));
  nor2   g430(.a(n464), .b(n453), .O(n489));
  nor2   g431(.a(n489), .b(n85), .O(n490));
  inv1   g432(.a(n489), .O(n491));
  nor2   g433(.a(n491), .b(G140), .O(n492));
  nor2   g434(.a(n492), .b(n490), .O(n493));
  inv1   g435(.a(n493), .O(G42));
  nor2   g436(.a(n426), .b(n420), .O(n495));
  inv1   g437(.a(n495), .O(n496));
  nor2   g438(.a(n446), .b(n434), .O(n497));
  inv1   g439(.a(n497), .O(n498));
  nor2   g440(.a(n498), .b(n496), .O(n499));
  inv1   g441(.a(n499), .O(n500));
  nor2   g442(.a(n353), .b(n338), .O(n501));
  inv1   g443(.a(n501), .O(n502));
  nor2   g444(.a(n373), .b(n363), .O(n503));
  inv1   g445(.a(n503), .O(n504));
  nor2   g446(.a(n504), .b(n502), .O(n505));
  inv1   g447(.a(n505), .O(n506));
  nor2   g448(.a(n506), .b(n500), .O(n507));
  inv1   g449(.a(n507), .O(n508));
  nor2   g450(.a(n473), .b(n467), .O(n509));
  inv1   g451(.a(n509), .O(n510));
  nor2   g452(.a(n489), .b(n483), .O(n511));
  inv1   g453(.a(n511), .O(n512));
  nor2   g454(.a(n512), .b(n510), .O(n513));
  inv1   g455(.a(n513), .O(n514));
  nor2   g456(.a(n399), .b(n389), .O(n515));
  inv1   g457(.a(n515), .O(n516));
  nor2   g458(.a(n454), .b(n407), .O(n517));
  inv1   g459(.a(n517), .O(n518));
  nor2   g460(.a(n518), .b(n516), .O(n519));
  inv1   g461(.a(n519), .O(n520));
  nor2   g462(.a(n520), .b(n514), .O(n521));
  inv1   g463(.a(n521), .O(n522));
  nor2   g464(.a(n522), .b(n508), .O(n523));
  inv1   g465(.a(n523), .O(n524));
  nor2   g466(.a(n323), .b(n321), .O(n525));
  inv1   g467(.a(n525), .O(n526));
  inv1   g468(.a(n218), .O(n527));
  nor2   g469(.a(n243), .b(n527), .O(n528));
  nor2   g470(.a(n528), .b(n346), .O(n529));
  nor2   g471(.a(n415), .b(n379), .O(n530));
  nor2   g472(.a(n530), .b(n529), .O(n531));
  nor2   g473(.a(n462), .b(n440), .O(n532));
  inv1   g474(.a(n532), .O(n533));
  nor2   g475(.a(n533), .b(n531), .O(n534));
  nor2   g476(.a(n534), .b(n442), .O(n535));
  nor2   g477(.a(n535), .b(n526), .O(n536));
  inv1   g478(.a(n170), .O(n537));
  nor2   g479(.a(n525), .b(n537), .O(n538));
  inv1   g480(.a(n323), .O(n539));
  nor2   g481(.a(n539), .b(n320), .O(n540));
  nor2   g482(.a(n395), .b(n460), .O(n541));
  inv1   g483(.a(n541), .O(n542));
  nor2   g484(.a(n542), .b(n441), .O(n543));
  inv1   g485(.a(n543), .O(n544));
  nor2   g486(.a(n544), .b(n540), .O(n545));
  inv1   g487(.a(n545), .O(n546));
  nor2   g488(.a(n546), .b(n538), .O(n547));
  nor2   g489(.a(n547), .b(n326), .O(n548));
  inv1   g490(.a(n548), .O(n549));
  nor2   g491(.a(n549), .b(n536), .O(n550));
  inv1   g492(.a(n550), .O(n551));
  nor2   g493(.a(n551), .b(n524), .O(n552));
  nor2   g494(.a(n462), .b(n321), .O(n553));
  inv1   g495(.a(n553), .O(n554));
  nor2   g496(.a(n554), .b(n441), .O(n555));
  nor2   g497(.a(G953), .b(G952), .O(n556));
  inv1   g498(.a(n556), .O(n557));
  nor2   g499(.a(n557), .b(n555), .O(n558));
  nor2   g500(.a(n558), .b(n552), .O(G75));
  nor2   g501(.a(n331), .b(n121), .O(n560));
  inv1   g502(.a(n560), .O(n561));
  nor2   g503(.a(n561), .b(n523), .O(n562));
  inv1   g504(.a(n562), .O(n563));
  nor2   g505(.a(n563), .b(n209), .O(n564));
  nor2   g506(.a(n328), .b(G952), .O(n565));
  nor2   g507(.a(n562), .b(n208), .O(n566));
  nor2   g508(.a(n566), .b(n565), .O(n567));
  inv1   g509(.a(n567), .O(n568));
  nor2   g510(.a(n568), .b(n564), .O(G51));
  nor2   g511(.a(n331), .b(n219), .O(n570));
  inv1   g512(.a(n570), .O(n571));
  nor2   g513(.a(n571), .b(n523), .O(n572));
  inv1   g514(.a(n572), .O(n573));
  nor2   g515(.a(n573), .b(n238), .O(n574));
  nor2   g516(.a(n572), .b(n237), .O(n575));
  nor2   g517(.a(n575), .b(n565), .O(n576));
  inv1   g518(.a(n576), .O(n577));
  nor2   g519(.a(n577), .b(n574), .O(G54));
  nor2   g520(.a(n331), .b(n285), .O(n579));
  inv1   g521(.a(n579), .O(n580));
  nor2   g522(.a(n580), .b(n523), .O(n581));
  nor2   g523(.a(n581), .b(n312), .O(n582));
  inv1   g524(.a(n581), .O(n583));
  nor2   g525(.a(n583), .b(n313), .O(n584));
  nor2   g526(.a(n584), .b(n565), .O(n585));
  inv1   g527(.a(n585), .O(n586));
  nor2   g528(.a(n586), .b(n582), .O(G60));
  nor2   g529(.a(n331), .b(n250), .O(n588));
  inv1   g530(.a(n588), .O(n589));
  nor2   g531(.a(n589), .b(n523), .O(n590));
  nor2   g532(.a(n590), .b(n277), .O(n591));
  inv1   g533(.a(n590), .O(n592));
  nor2   g534(.a(n592), .b(n278), .O(n593));
  nor2   g535(.a(n593), .b(n565), .O(n594));
  inv1   g536(.a(n594), .O(n595));
  nor2   g537(.a(n595), .b(n591), .O(G63));
  nor2   g538(.a(n331), .b(n101), .O(n597));
  inv1   g539(.a(n597), .O(n598));
  nor2   g540(.a(n598), .b(n523), .O(n599));
  inv1   g541(.a(n599), .O(n600));
  nor2   g542(.a(n600), .b(n99), .O(n601));
  inv1   g543(.a(n99), .O(n602));
  nor2   g544(.a(n599), .b(n602), .O(n603));
  nor2   g545(.a(n603), .b(n565), .O(n604));
  inv1   g546(.a(n604), .O(n605));
  nor2   g547(.a(n605), .b(n601), .O(G66));
  nor2   g548(.a(n507), .b(G953), .O(n607));
  nor2   g549(.a(n328), .b(G224), .O(n608));
  nor2   g550(.a(n608), .b(n607), .O(n609));
  nor2   g551(.a(n609), .b(n193), .O(n610));
  inv1   g552(.a(n609), .O(n611));
  nor2   g553(.a(n611), .b(n194), .O(n612));
  nor2   g554(.a(n612), .b(n610), .O(n613));
  nor2   g555(.a(n613), .b(n329), .O(n614));
  inv1   g556(.a(n614), .O(G69));
  nor2   g557(.a(n521), .b(G953), .O(n616));
  nor2   g558(.a(n328), .b(G227), .O(n617));
  nor2   g559(.a(n617), .b(n383), .O(n618));
  inv1   g560(.a(n618), .O(n619));
  nor2   g561(.a(n619), .b(n616), .O(n620));
  nor2   g562(.a(n151), .b(n89), .O(n621));
  nor2   g563(.a(n153), .b(n87), .O(n622));
  nor2   g564(.a(n622), .b(n621), .O(n623));
  nor2   g565(.a(n623), .b(n383), .O(n624));
  inv1   g566(.a(n624), .O(n625));
  nor2   g567(.a(n625), .b(n620), .O(n626));
  inv1   g568(.a(n620), .O(n627));
  nor2   g569(.a(n624), .b(n627), .O(n628));
  nor2   g570(.a(n628), .b(n626), .O(G72));
  nor2   g571(.a(n331), .b(n110), .O(n630));
  inv1   g572(.a(n630), .O(n631));
  nor2   g573(.a(n631), .b(n523), .O(n632));
  inv1   g574(.a(n632), .O(n633));
  nor2   g575(.a(n633), .b(n160), .O(n634));
  nor2   g576(.a(n632), .b(n159), .O(n635));
  nor2   g577(.a(n635), .b(n565), .O(n636));
  inv1   g578(.a(n636), .O(n637));
  nor2   g579(.a(n637), .b(n634), .O(G57));
endmodule


