// Benchmark "c7552_blif" written by ABC on Sun Mar 24 18:35:07 2019

module c7552_blif  ( 
    G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47,
    G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65,
    G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83,
    G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110,
    G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133, G134,
    G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, G155, G156,
    G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, G167, G168,
    G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179, G180,
    G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G216,
    G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227, G228,
    G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239, G240,
    ING339 , G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492,
    G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247,
    G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737,
    G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427,
    G4432, G4437, G4526, G4528,
    G339, G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492,
    G490, G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552,
    G550, G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526,
    G524, G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446,
    G284, G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264,
    G270, G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416,
    G249, G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333,
    G336, G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471,
    G359, G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399  );
  input  G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41,
    G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63,
    G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81,
    G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106,
    G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130,
    G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154,
    G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166,
    G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190,
    G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202,
    G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214,
    G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226,
    G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238,
    G239, G240, ING339 , G1197, G1455, G1459, G1462, G1469, G1480, G1486,
    G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239,
    G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729,
    G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420,
    G4427, G4432, G4437, G4526, G4528;
  output G339, G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492,
    G490, G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552,
    G550, G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526,
    G524, G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446,
    G284, G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264,
    G270, G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416,
    G249, G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333,
    G336, G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471,
    G359, G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399;
  wire n317, n319, n320, n321, n322, n323, n324, n325, n326, n327, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n339, n340, n341, n342,
    n343, n344, n345, n346, n347, n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n359, n360, n362, n363, n364, n365, n366, n368, n369, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
    n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
    n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
    n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
    n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
    n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
    n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
    n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
    n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
    n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
    n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
    n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
    n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
    n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
    n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
    n1389, n1390, n1391, n1392, n1393, n1394, n1396, n1397, n1399, n1400,
    n1401, n1402, n1403, n1404, n1406, n1407, n1409, n1410, n1411, n1412,
    n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1421, n1422, n1424,
    n1425, n1426, n1427, n1429, n1430, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
    n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
    n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
    n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1605, n1606, n1607,
    n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
    n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
    n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
    n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
    n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
    n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
    n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
    n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
    n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
    n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
    n1939, n1940, n1941, n1942, n1943, n1945, n1946, n1947, n1949, n1950,
    n1951, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1974,
    n1975, n1976, n1977, n1978, n1979, n1981, n1982, n1984, n1985, n1986,
    n1987, n1988, n1989, n1990, n1991, n1993, n1994, n1995, n1996, n1997,
    n1998, n2000, n2001, n2002, n2004, n2005, n2006, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2020, n2021,
    n2022, n2023, n2024, n2025, n2027, n2028, n2029, n2030, n2031, n2032,
    n2033, n2034, n2035, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2049, n2050, n2052, n2053, n2054, n2055,
    n2056, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
    n2067, n2068, n2070, n2071, n2072, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2088, n2089,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2099, n2100, n2101,
    n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2112, n2113,
    n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2122, n2123, n2124,
    n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2134, n2135,
    n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
    n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
    n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
    n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
    n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
    n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2223, n2224, n2225, n2226, n2227,
    n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
    n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
    n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
    n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
    n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
    n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
    n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
    n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
    n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
    n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
    n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
    n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
    n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
    n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
    n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
    n2480, n2481;
  inv1   g0000(.a(G15), .O(G279));
  nor2   g0001(.a(G57), .b(G5), .O(n317));
  inv1   g0002(.a(n317), .O(G402));
  inv1   g0003(.a(G150), .O(n319));
  inv1   g0004(.a(G184), .O(n320));
  nor2   g0005(.a(n320), .b(n319), .O(n321));
  inv1   g0006(.a(n321), .O(n322));
  inv1   g0007(.a(G228), .O(n323));
  inv1   g0008(.a(G240), .O(n324));
  nor2   g0009(.a(n324), .b(n323), .O(n325));
  inv1   g0010(.a(n325), .O(n326));
  nor2   g0011(.a(n326), .b(n322), .O(n327));
  inv1   g0012(.a(n327), .O(G404));
  inv1   g0013(.a(G152), .O(n329));
  inv1   g0014(.a(G210), .O(n330));
  nor2   g0015(.a(n330), .b(n329), .O(n331));
  inv1   g0016(.a(n331), .O(n332));
  inv1   g0017(.a(G218), .O(n333));
  inv1   g0018(.a(G230), .O(n334));
  nor2   g0019(.a(n334), .b(n333), .O(n335));
  inv1   g0020(.a(n335), .O(n336));
  nor2   g0021(.a(n336), .b(n332), .O(n337));
  inv1   g0022(.a(n337), .O(G406));
  inv1   g0023(.a(G182), .O(n339));
  inv1   g0024(.a(G183), .O(n340));
  nor2   g0025(.a(n340), .b(n339), .O(n341));
  inv1   g0026(.a(n341), .O(n342));
  inv1   g0027(.a(G185), .O(n343));
  inv1   g0028(.a(G186), .O(n344));
  nor2   g0029(.a(n344), .b(n343), .O(n345));
  inv1   g0030(.a(n345), .O(n346));
  nor2   g0031(.a(n346), .b(n342), .O(n347));
  inv1   g0032(.a(n347), .O(G408));
  inv1   g0033(.a(G162), .O(n349));
  inv1   g0034(.a(G172), .O(n350));
  nor2   g0035(.a(n350), .b(n349), .O(n351));
  inv1   g0036(.a(n351), .O(n352));
  inv1   g0037(.a(G188), .O(n353));
  inv1   g0038(.a(G199), .O(n354));
  nor2   g0039(.a(n354), .b(n353), .O(n355));
  inv1   g0040(.a(n355), .O(n356));
  nor2   g0041(.a(n356), .b(n352), .O(n357));
  inv1   g0042(.a(n357), .O(G410));
  inv1   g0043(.a(G1197), .O(n359));
  nor2   g0044(.a(n359), .b(G5), .O(n360));
  inv1   g0045(.a(n360), .O(G284));
  inv1   g0046(.a(G134), .O(n362));
  inv1   g0047(.a(G133), .O(n363));
  nor2   g0048(.a(n363), .b(G5), .O(n364));
  inv1   g0049(.a(n364), .O(n365));
  nor2   g0050(.a(n365), .b(n362), .O(n366));
  inv1   g0051(.a(n366), .O(G292));
  inv1   g0052(.a(G1), .O(n368));
  inv1   g0053(.a(G163), .O(n369));
  nor2   g0054(.a(n369), .b(n368), .O(G278));
  inv1   g0055(.a(G4526), .O(n371));
  inv1   g0056(.a(G41), .O(n372));
  nor2   g0057(.a(n372), .b(G18), .O(n373));
  inv1   g0058(.a(n373), .O(n374));
  nor2   g0059(.a(n374), .b(G3701), .O(n375));
  inv1   g0060(.a(G3701), .O(n376));
  nor2   g0061(.a(G41), .b(G18), .O(n377));
  inv1   g0062(.a(n377), .O(n378));
  nor2   g0063(.a(n378), .b(n376), .O(n379));
  nor2   g0064(.a(n379), .b(n375), .O(n380));
  inv1   g0065(.a(n380), .O(n381));
  nor2   g0066(.a(n381), .b(n371), .O(n382));
  nor2   g0067(.a(n380), .b(G4526), .O(n383));
  nor2   g0068(.a(n383), .b(n382), .O(G373));
  inv1   g0069(.a(G1496), .O(n385));
  inv1   g0070(.a(G4528), .O(n386));
  nor2   g0071(.a(n386), .b(n385), .O(n387));
  inv1   g0072(.a(G1492), .O(n388));
  nor2   g0073(.a(n386), .b(n388), .O(n389));
  nor2   g0074(.a(n389), .b(G38), .O(n390));
  inv1   g0075(.a(n390), .O(n391));
  nor2   g0076(.a(n391), .b(n387), .O(n392));
  inv1   g0077(.a(n392), .O(n393));
  inv1   g0078(.a(G9), .O(n394));
  inv1   g0079(.a(G12), .O(n395));
  nor2   g0080(.a(n395), .b(n394), .O(n396));
  inv1   g0081(.a(G18), .O(n397));
  nor2   g0082(.a(G153), .b(n397), .O(n398));
  nor2   g0083(.a(n398), .b(n396), .O(n399));
  inv1   g0084(.a(n399), .O(n400));
  nor2   g0085(.a(n400), .b(G2256), .O(n401));
  inv1   g0086(.a(G2256), .O(n402));
  nor2   g0087(.a(n399), .b(n402), .O(n403));
  nor2   g0088(.a(n403), .b(n401), .O(n404));
  inv1   g0089(.a(n404), .O(n405));
  inv1   g0090(.a(G2253), .O(n406));
  nor2   g0091(.a(G154), .b(n397), .O(n407));
  nor2   g0092(.a(n407), .b(n396), .O(n408));
  nor2   g0093(.a(n408), .b(n406), .O(n409));
  nor2   g0094(.a(G155), .b(n397), .O(n410));
  nor2   g0095(.a(n410), .b(n396), .O(n411));
  inv1   g0096(.a(n411), .O(n412));
  nor2   g0097(.a(n412), .b(G2247), .O(n413));
  inv1   g0098(.a(G2247), .O(n414));
  nor2   g0099(.a(n411), .b(n414), .O(n415));
  nor2   g0100(.a(n415), .b(n413), .O(n416));
  inv1   g0101(.a(n416), .O(n417));
  nor2   g0102(.a(G156), .b(n397), .O(n418));
  nor2   g0103(.a(n418), .b(n396), .O(n419));
  inv1   g0104(.a(n419), .O(n420));
  nor2   g0105(.a(n420), .b(G2239), .O(n421));
  inv1   g0106(.a(n421), .O(n422));
  nor2   g0107(.a(n422), .b(n417), .O(n423));
  nor2   g0108(.a(n423), .b(n413), .O(n424));
  inv1   g0109(.a(n424), .O(n425));
  nor2   g0110(.a(n425), .b(n409), .O(n426));
  inv1   g0111(.a(n426), .O(n427));
  inv1   g0112(.a(n408), .O(n428));
  nor2   g0113(.a(n428), .b(G2253), .O(n429));
  inv1   g0114(.a(G2239), .O(n430));
  nor2   g0115(.a(n419), .b(n430), .O(n431));
  nor2   g0116(.a(n431), .b(n417), .O(n432));
  nor2   g0117(.a(n432), .b(n413), .O(n433));
  nor2   g0118(.a(n433), .b(n429), .O(n434));
  inv1   g0119(.a(n434), .O(n435));
  nor2   g0120(.a(n435), .b(n427), .O(n436));
  inv1   g0121(.a(n436), .O(n437));
  nor2   g0122(.a(n437), .b(n405), .O(n438));
  inv1   g0123(.a(n438), .O(n439));
  inv1   g0124(.a(G234), .O(n440));
  nor2   g0125(.a(n440), .b(n397), .O(n441));
  inv1   g0126(.a(G130), .O(n442));
  nor2   g0127(.a(n442), .b(G18), .O(n443));
  nor2   g0128(.a(n443), .b(n441), .O(n444));
  nor2   g0129(.a(n444), .b(G3729), .O(n445));
  inv1   g0130(.a(G3729), .O(n446));
  inv1   g0131(.a(n444), .O(n447));
  nor2   g0132(.a(n447), .b(n446), .O(n448));
  nor2   g0133(.a(n448), .b(n445), .O(n449));
  inv1   g0134(.a(n449), .O(n450));
  inv1   g0135(.a(G233), .O(n451));
  nor2   g0136(.a(n451), .b(n397), .O(n452));
  inv1   g0137(.a(G127), .O(n453));
  nor2   g0138(.a(n453), .b(G18), .O(n454));
  nor2   g0139(.a(n454), .b(n452), .O(n455));
  nor2   g0140(.a(n455), .b(G3737), .O(n456));
  inv1   g0141(.a(G3737), .O(n457));
  inv1   g0142(.a(n455), .O(n458));
  nor2   g0143(.a(n458), .b(n457), .O(n459));
  nor2   g0144(.a(n459), .b(n456), .O(n460));
  inv1   g0145(.a(n460), .O(n461));
  nor2   g0146(.a(n461), .b(n450), .O(n462));
  inv1   g0147(.a(n462), .O(n463));
  inv1   g0148(.a(G231), .O(n464));
  nor2   g0149(.a(n464), .b(n397), .O(n465));
  inv1   g0150(.a(G100), .O(n466));
  nor2   g0151(.a(n466), .b(G18), .O(n467));
  nor2   g0152(.a(n467), .b(n465), .O(n468));
  nor2   g0153(.a(n468), .b(G3749), .O(n469));
  inv1   g0154(.a(G3749), .O(n470));
  inv1   g0155(.a(n468), .O(n471));
  nor2   g0156(.a(n471), .b(n470), .O(n472));
  nor2   g0157(.a(n472), .b(n469), .O(n473));
  inv1   g0158(.a(n473), .O(n474));
  inv1   g0159(.a(G232), .O(n475));
  nor2   g0160(.a(n475), .b(n397), .O(n476));
  inv1   g0161(.a(G124), .O(n477));
  nor2   g0162(.a(n477), .b(G18), .O(n478));
  nor2   g0163(.a(n478), .b(n476), .O(n479));
  nor2   g0164(.a(n479), .b(G3743), .O(n480));
  inv1   g0165(.a(G3743), .O(n481));
  inv1   g0166(.a(n479), .O(n482));
  nor2   g0167(.a(n482), .b(n481), .O(n483));
  nor2   g0168(.a(n483), .b(n480), .O(n484));
  inv1   g0169(.a(n484), .O(n485));
  nor2   g0170(.a(n485), .b(n474), .O(n486));
  inv1   g0171(.a(n486), .O(n487));
  nor2   g0172(.a(n487), .b(n463), .O(n488));
  inv1   g0173(.a(n488), .O(n489));
  inv1   g0174(.a(G235), .O(n490));
  nor2   g0175(.a(n490), .b(n397), .O(n491));
  inv1   g0176(.a(G103), .O(n492));
  nor2   g0177(.a(n492), .b(G18), .O(n493));
  nor2   g0178(.a(n493), .b(n491), .O(n494));
  nor2   g0179(.a(n494), .b(G3723), .O(n495));
  inv1   g0180(.a(G3723), .O(n496));
  inv1   g0181(.a(n494), .O(n497));
  nor2   g0182(.a(n497), .b(n496), .O(n498));
  nor2   g0183(.a(n498), .b(n495), .O(n499));
  inv1   g0184(.a(n499), .O(n500));
  inv1   g0185(.a(G236), .O(n501));
  nor2   g0186(.a(n501), .b(n397), .O(n502));
  inv1   g0187(.a(G23), .O(n503));
  nor2   g0188(.a(n503), .b(G18), .O(n504));
  nor2   g0189(.a(n504), .b(n502), .O(n505));
  nor2   g0190(.a(n505), .b(G3717), .O(n506));
  inv1   g0191(.a(G3717), .O(n507));
  inv1   g0192(.a(n505), .O(n508));
  nor2   g0193(.a(n508), .b(n507), .O(n509));
  nor2   g0194(.a(n509), .b(n506), .O(n510));
  inv1   g0195(.a(n510), .O(n511));
  nor2   g0196(.a(n511), .b(n500), .O(n512));
  inv1   g0197(.a(n512), .O(n513));
  inv1   g0198(.a(G3711), .O(n514));
  inv1   g0199(.a(G237), .O(n515));
  nor2   g0200(.a(n515), .b(n397), .O(n516));
  inv1   g0201(.a(G26), .O(n517));
  nor2   g0202(.a(n517), .b(G18), .O(n518));
  nor2   g0203(.a(n518), .b(n516), .O(n519));
  inv1   g0204(.a(n519), .O(n520));
  nor2   g0205(.a(n520), .b(n514), .O(n521));
  nor2   g0206(.a(n519), .b(G3711), .O(n522));
  inv1   g0207(.a(G3705), .O(n523));
  inv1   g0208(.a(G238), .O(n524));
  nor2   g0209(.a(n524), .b(n397), .O(n525));
  inv1   g0210(.a(G29), .O(n526));
  nor2   g0211(.a(n526), .b(G18), .O(n527));
  nor2   g0212(.a(n527), .b(n525), .O(n528));
  inv1   g0213(.a(n528), .O(n529));
  nor2   g0214(.a(n529), .b(n523), .O(n530));
  nor2   g0215(.a(n528), .b(G3705), .O(n531));
  nor2   g0216(.a(n531), .b(n375), .O(n532));
  nor2   g0217(.a(n532), .b(n530), .O(n533));
  nor2   g0218(.a(n533), .b(n522), .O(n534));
  nor2   g0219(.a(n534), .b(n521), .O(n535));
  inv1   g0220(.a(n535), .O(n536));
  nor2   g0221(.a(n536), .b(n513), .O(n537));
  nor2   g0222(.a(n506), .b(n495), .O(n538));
  nor2   g0223(.a(n538), .b(n498), .O(n539));
  nor2   g0224(.a(n539), .b(n537), .O(n540));
  nor2   g0225(.a(n540), .b(n489), .O(n541));
  inv1   g0226(.a(n445), .O(n542));
  nor2   g0227(.a(n461), .b(n542), .O(n543));
  nor2   g0228(.a(n543), .b(n456), .O(n544));
  nor2   g0229(.a(n544), .b(n483), .O(n545));
  nor2   g0230(.a(n545), .b(n480), .O(n546));
  nor2   g0231(.a(n546), .b(n472), .O(n547));
  nor2   g0232(.a(n547), .b(n469), .O(n548));
  inv1   g0233(.a(n548), .O(n549));
  nor2   g0234(.a(n549), .b(n541), .O(n550));
  inv1   g0235(.a(G219), .O(n551));
  nor2   g0236(.a(n551), .b(n397), .O(n552));
  inv1   g0237(.a(G66), .O(n553));
  nor2   g0238(.a(n553), .b(G18), .O(n554));
  nor2   g0239(.a(n554), .b(n552), .O(n555));
  nor2   g0240(.a(n555), .b(G4437), .O(n556));
  inv1   g0241(.a(G4437), .O(n557));
  inv1   g0242(.a(n555), .O(n558));
  nor2   g0243(.a(n558), .b(n557), .O(n559));
  nor2   g0244(.a(n559), .b(n556), .O(n560));
  inv1   g0245(.a(n560), .O(n561));
  inv1   g0246(.a(G4432), .O(n562));
  inv1   g0247(.a(G220), .O(n563));
  nor2   g0248(.a(n563), .b(n397), .O(n564));
  inv1   g0249(.a(G50), .O(n565));
  nor2   g0250(.a(n565), .b(G18), .O(n566));
  nor2   g0251(.a(n566), .b(n564), .O(n567));
  inv1   g0252(.a(n567), .O(n568));
  nor2   g0253(.a(n568), .b(n562), .O(n569));
  inv1   g0254(.a(G221), .O(n570));
  nor2   g0255(.a(n570), .b(n397), .O(n571));
  inv1   g0256(.a(G32), .O(n572));
  nor2   g0257(.a(n572), .b(G18), .O(n573));
  nor2   g0258(.a(n573), .b(n571), .O(n574));
  nor2   g0259(.a(n574), .b(G4427), .O(n575));
  inv1   g0260(.a(G4427), .O(n576));
  inv1   g0261(.a(n574), .O(n577));
  nor2   g0262(.a(n577), .b(n576), .O(n578));
  nor2   g0263(.a(n578), .b(n575), .O(n579));
  inv1   g0264(.a(n579), .O(n580));
  inv1   g0265(.a(G222), .O(n581));
  nor2   g0266(.a(n581), .b(n397), .O(n582));
  inv1   g0267(.a(G35), .O(n583));
  nor2   g0268(.a(n583), .b(G18), .O(n584));
  nor2   g0269(.a(n584), .b(n582), .O(n585));
  nor2   g0270(.a(n585), .b(G4420), .O(n586));
  inv1   g0271(.a(n586), .O(n587));
  nor2   g0272(.a(n587), .b(n580), .O(n588));
  nor2   g0273(.a(n588), .b(n575), .O(n589));
  inv1   g0274(.a(n589), .O(n590));
  nor2   g0275(.a(n590), .b(n569), .O(n591));
  inv1   g0276(.a(n591), .O(n592));
  nor2   g0277(.a(n567), .b(G4432), .O(n593));
  inv1   g0278(.a(G4420), .O(n594));
  inv1   g0279(.a(n585), .O(n595));
  nor2   g0280(.a(n595), .b(n594), .O(n596));
  nor2   g0281(.a(n596), .b(n580), .O(n597));
  nor2   g0282(.a(n597), .b(n575), .O(n598));
  nor2   g0283(.a(n598), .b(n593), .O(n599));
  inv1   g0284(.a(n599), .O(n600));
  nor2   g0285(.a(n600), .b(n592), .O(n601));
  inv1   g0286(.a(n601), .O(n602));
  nor2   g0287(.a(n602), .b(n561), .O(n603));
  inv1   g0288(.a(n603), .O(n604));
  inv1   g0289(.a(G223), .O(n605));
  nor2   g0290(.a(n605), .b(n397), .O(n606));
  inv1   g0291(.a(G47), .O(n607));
  nor2   g0292(.a(n607), .b(G18), .O(n608));
  nor2   g0293(.a(n608), .b(n606), .O(n609));
  nor2   g0294(.a(n609), .b(G4415), .O(n610));
  inv1   g0295(.a(G4415), .O(n611));
  inv1   g0296(.a(n609), .O(n612));
  nor2   g0297(.a(n612), .b(n611), .O(n613));
  nor2   g0298(.a(n613), .b(n610), .O(n614));
  inv1   g0299(.a(n614), .O(n615));
  inv1   g0300(.a(G224), .O(n616));
  nor2   g0301(.a(n616), .b(n397), .O(n617));
  inv1   g0302(.a(G121), .O(n618));
  nor2   g0303(.a(n618), .b(G18), .O(n619));
  nor2   g0304(.a(n619), .b(n617), .O(n620));
  nor2   g0305(.a(n620), .b(G4410), .O(n621));
  inv1   g0306(.a(G4410), .O(n622));
  inv1   g0307(.a(n620), .O(n623));
  nor2   g0308(.a(n623), .b(n622), .O(n624));
  nor2   g0309(.a(n624), .b(n621), .O(n625));
  inv1   g0310(.a(n625), .O(n626));
  nor2   g0311(.a(n626), .b(n615), .O(n627));
  inv1   g0312(.a(n627), .O(n628));
  inv1   g0313(.a(G226), .O(n629));
  nor2   g0314(.a(n629), .b(n397), .O(n630));
  inv1   g0315(.a(G97), .O(n631));
  nor2   g0316(.a(n631), .b(G18), .O(n632));
  nor2   g0317(.a(n632), .b(n630), .O(n633));
  nor2   g0318(.a(n633), .b(G4400), .O(n634));
  inv1   g0319(.a(G4400), .O(n635));
  inv1   g0320(.a(n633), .O(n636));
  nor2   g0321(.a(n636), .b(n635), .O(n637));
  nor2   g0322(.a(n637), .b(n634), .O(n638));
  inv1   g0323(.a(n638), .O(n639));
  inv1   g0324(.a(G217), .O(n640));
  nor2   g0325(.a(n640), .b(n397), .O(n641));
  inv1   g0326(.a(G118), .O(n642));
  nor2   g0327(.a(n642), .b(G18), .O(n643));
  nor2   g0328(.a(n643), .b(n641), .O(n644));
  nor2   g0329(.a(n644), .b(G4394), .O(n645));
  inv1   g0330(.a(G4394), .O(n646));
  inv1   g0331(.a(n644), .O(n647));
  nor2   g0332(.a(n647), .b(n646), .O(n648));
  nor2   g0333(.a(n648), .b(n645), .O(n649));
  inv1   g0334(.a(n649), .O(n650));
  nor2   g0335(.a(n650), .b(n639), .O(n651));
  inv1   g0336(.a(n651), .O(n652));
  inv1   g0337(.a(G225), .O(n653));
  nor2   g0338(.a(n653), .b(n397), .O(n654));
  inv1   g0339(.a(G94), .O(n655));
  nor2   g0340(.a(n655), .b(G18), .O(n656));
  nor2   g0341(.a(n656), .b(n654), .O(n657));
  nor2   g0342(.a(n657), .b(G4405), .O(n658));
  inv1   g0343(.a(G4405), .O(n659));
  inv1   g0344(.a(n657), .O(n660));
  nor2   g0345(.a(n660), .b(n659), .O(n661));
  nor2   g0346(.a(n661), .b(n658), .O(n662));
  inv1   g0347(.a(n662), .O(n663));
  nor2   g0348(.a(n663), .b(n652), .O(n664));
  inv1   g0349(.a(n664), .O(n665));
  nor2   g0350(.a(n665), .b(n628), .O(n666));
  inv1   g0351(.a(n666), .O(n667));
  nor2   g0352(.a(n667), .b(n604), .O(n668));
  inv1   g0353(.a(n668), .O(n669));
  nor2   g0354(.a(n669), .b(n550), .O(n670));
  inv1   g0355(.a(n645), .O(n671));
  nor2   g0356(.a(n671), .b(n639), .O(n672));
  inv1   g0357(.a(n672), .O(n673));
  nor2   g0358(.a(n673), .b(n661), .O(n674));
  nor2   g0359(.a(n674), .b(n658), .O(n675));
  nor2   g0360(.a(n675), .b(n628), .O(n676));
  inv1   g0361(.a(n634), .O(n677));
  nor2   g0362(.a(n663), .b(n677), .O(n678));
  inv1   g0363(.a(n678), .O(n679));
  nor2   g0364(.a(n679), .b(n628), .O(n680));
  inv1   g0365(.a(n621), .O(n681));
  nor2   g0366(.a(n681), .b(n613), .O(n682));
  nor2   g0367(.a(n682), .b(n610), .O(n683));
  inv1   g0368(.a(n683), .O(n684));
  nor2   g0369(.a(n684), .b(n680), .O(n685));
  inv1   g0370(.a(n685), .O(n686));
  nor2   g0371(.a(n686), .b(n676), .O(n687));
  inv1   g0372(.a(n687), .O(n688));
  nor2   g0373(.a(n531), .b(n530), .O(n689));
  inv1   g0374(.a(n689), .O(n690));
  nor2   g0375(.a(n690), .b(n381), .O(n691));
  inv1   g0376(.a(n691), .O(n692));
  nor2   g0377(.a(n522), .b(n521), .O(n693));
  inv1   g0378(.a(n693), .O(n694));
  nor2   g0379(.a(n694), .b(n371), .O(n695));
  inv1   g0380(.a(n695), .O(n696));
  nor2   g0381(.a(n696), .b(n692), .O(n697));
  inv1   g0382(.a(n697), .O(n698));
  nor2   g0383(.a(n698), .b(n513), .O(n699));
  inv1   g0384(.a(n699), .O(n700));
  nor2   g0385(.a(n667), .b(n489), .O(n701));
  inv1   g0386(.a(n701), .O(n702));
  nor2   g0387(.a(n702), .b(n700), .O(n703));
  nor2   g0388(.a(n703), .b(n688), .O(n704));
  nor2   g0389(.a(n704), .b(n604), .O(n705));
  nor2   g0390(.a(n589), .b(n569), .O(n706));
  nor2   g0391(.a(n706), .b(n593), .O(n707));
  inv1   g0392(.a(n707), .O(n708));
  nor2   g0393(.a(n708), .b(n556), .O(n709));
  nor2   g0394(.a(n709), .b(n559), .O(n710));
  nor2   g0395(.a(n710), .b(n705), .O(n711));
  inv1   g0396(.a(n711), .O(n712));
  nor2   g0397(.a(n712), .b(n670), .O(n713));
  inv1   g0398(.a(G135), .O(n714));
  nor2   g0399(.a(n714), .b(G18), .O(n715));
  inv1   g0400(.a(G158), .O(n716));
  nor2   g0401(.a(n716), .b(n397), .O(n717));
  nor2   g0402(.a(n717), .b(n715), .O(n718));
  nor2   g0403(.a(n718), .b(G2230), .O(n719));
  inv1   g0404(.a(G2230), .O(n720));
  inv1   g0405(.a(n718), .O(n721));
  nor2   g0406(.a(n721), .b(n720), .O(n722));
  nor2   g0407(.a(n722), .b(n719), .O(n723));
  inv1   g0408(.a(n723), .O(n724));
  inv1   g0409(.a(G144), .O(n725));
  nor2   g0410(.a(n725), .b(G18), .O(n726));
  inv1   g0411(.a(G159), .O(n727));
  nor2   g0412(.a(n727), .b(n397), .O(n728));
  nor2   g0413(.a(n728), .b(n726), .O(n729));
  nor2   g0414(.a(n729), .b(G2224), .O(n730));
  inv1   g0415(.a(G2224), .O(n731));
  inv1   g0416(.a(n729), .O(n732));
  nor2   g0417(.a(n732), .b(n731), .O(n733));
  nor2   g0418(.a(n733), .b(n730), .O(n734));
  inv1   g0419(.a(n734), .O(n735));
  nor2   g0420(.a(n735), .b(n724), .O(n736));
  inv1   g0421(.a(n736), .O(n737));
  inv1   g0422(.a(G138), .O(n738));
  nor2   g0423(.a(n738), .b(G18), .O(n739));
  inv1   g0424(.a(G160), .O(n740));
  nor2   g0425(.a(n740), .b(n397), .O(n741));
  nor2   g0426(.a(n741), .b(n739), .O(n742));
  nor2   g0427(.a(n742), .b(G2218), .O(n743));
  inv1   g0428(.a(G2218), .O(n744));
  inv1   g0429(.a(n742), .O(n745));
  nor2   g0430(.a(n745), .b(n744), .O(n746));
  nor2   g0431(.a(n746), .b(n743), .O(n747));
  inv1   g0432(.a(n747), .O(n748));
  inv1   g0433(.a(G147), .O(n749));
  nor2   g0434(.a(n749), .b(G18), .O(n750));
  inv1   g0435(.a(G151), .O(n751));
  nor2   g0436(.a(n751), .b(n397), .O(n752));
  nor2   g0437(.a(n752), .b(n750), .O(n753));
  nor2   g0438(.a(n753), .b(G2211), .O(n754));
  inv1   g0439(.a(G2211), .O(n755));
  inv1   g0440(.a(n753), .O(n756));
  nor2   g0441(.a(n756), .b(n755), .O(n757));
  nor2   g0442(.a(n757), .b(n754), .O(n758));
  inv1   g0443(.a(n758), .O(n759));
  nor2   g0444(.a(n759), .b(n748), .O(n760));
  inv1   g0445(.a(n760), .O(n761));
  nor2   g0446(.a(n761), .b(n737), .O(n762));
  inv1   g0447(.a(n762), .O(n763));
  nor2   g0448(.a(G157), .b(n397), .O(n764));
  nor2   g0449(.a(n764), .b(n396), .O(n765));
  inv1   g0450(.a(n765), .O(n766));
  nor2   g0451(.a(n766), .b(G2236), .O(n767));
  inv1   g0452(.a(G2236), .O(n768));
  nor2   g0453(.a(n765), .b(n768), .O(n769));
  nor2   g0454(.a(n769), .b(n767), .O(n770));
  inv1   g0455(.a(n770), .O(n771));
  nor2   g0456(.a(n771), .b(n763), .O(n772));
  inv1   g0457(.a(n772), .O(n773));
  nor2   g0458(.a(n773), .b(n713), .O(n774));
  inv1   g0459(.a(n774), .O(n775));
  nor2   g0460(.a(n775), .b(n439), .O(n776));
  inv1   g0461(.a(n754), .O(n777));
  nor2   g0462(.a(n777), .b(n748), .O(n778));
  nor2   g0463(.a(n778), .b(n743), .O(n779));
  nor2   g0464(.a(n779), .b(n733), .O(n780));
  nor2   g0465(.a(n780), .b(n730), .O(n781));
  nor2   g0466(.a(n781), .b(n722), .O(n782));
  nor2   g0467(.a(n782), .b(n719), .O(n783));
  inv1   g0468(.a(n783), .O(n784));
  nor2   g0469(.a(n784), .b(n767), .O(n785));
  nor2   g0470(.a(n785), .b(n769), .O(n786));
  inv1   g0471(.a(n786), .O(n787));
  nor2   g0472(.a(n787), .b(n439), .O(n788));
  nor2   g0473(.a(n429), .b(n425), .O(n789));
  nor2   g0474(.a(n789), .b(n409), .O(n790));
  inv1   g0475(.a(n790), .O(n791));
  nor2   g0476(.a(n791), .b(n403), .O(n792));
  nor2   g0477(.a(n792), .b(n401), .O(n793));
  inv1   g0478(.a(n793), .O(n794));
  nor2   g0479(.a(n794), .b(n788), .O(n795));
  inv1   g0480(.a(n795), .O(n796));
  nor2   g0481(.a(n796), .b(n776), .O(n797));
  nor2   g0482(.a(G216), .b(n397), .O(n798));
  nor2   g0483(.a(n798), .b(n396), .O(n799));
  inv1   g0484(.a(n799), .O(n800));
  nor2   g0485(.a(n800), .b(G1469), .O(n801));
  inv1   g0486(.a(G1469), .O(n802));
  nor2   g0487(.a(n799), .b(n802), .O(n803));
  nor2   g0488(.a(n803), .b(n801), .O(n804));
  inv1   g0489(.a(n804), .O(n805));
  nor2   g0490(.a(G209), .b(n397), .O(n806));
  nor2   g0491(.a(n806), .b(n396), .O(n807));
  inv1   g0492(.a(n807), .O(n808));
  nor2   g0493(.a(n808), .b(G1462), .O(n809));
  inv1   g0494(.a(G1462), .O(n810));
  nor2   g0495(.a(n807), .b(n810), .O(n811));
  nor2   g0496(.a(n811), .b(n809), .O(n812));
  inv1   g0497(.a(n812), .O(n813));
  nor2   g0498(.a(n813), .b(n805), .O(n814));
  inv1   g0499(.a(n814), .O(n815));
  nor2   g0500(.a(G214), .b(n397), .O(n816));
  nor2   g0501(.a(n816), .b(n396), .O(n817));
  inv1   g0502(.a(n817), .O(n818));
  nor2   g0503(.a(n818), .b(G1480), .O(n819));
  inv1   g0504(.a(G1480), .O(n820));
  nor2   g0505(.a(n817), .b(n820), .O(n821));
  nor2   g0506(.a(n821), .b(n819), .O(n822));
  inv1   g0507(.a(n822), .O(n823));
  nor2   g0508(.a(G215), .b(n397), .O(n824));
  nor2   g0509(.a(n824), .b(n396), .O(n825));
  inv1   g0510(.a(n825), .O(n826));
  nor2   g0511(.a(n826), .b(G106), .O(n827));
  inv1   g0512(.a(G106), .O(n828));
  nor2   g0513(.a(n825), .b(n828), .O(n829));
  nor2   g0514(.a(n829), .b(n827), .O(n830));
  inv1   g0515(.a(n830), .O(n831));
  nor2   g0516(.a(n831), .b(n823), .O(n832));
  inv1   g0517(.a(n832), .O(n833));
  nor2   g0518(.a(n833), .b(n815), .O(n834));
  inv1   g0519(.a(n834), .O(n835));
  nor2   g0520(.a(G213), .b(n397), .O(n836));
  nor2   g0521(.a(n836), .b(n396), .O(n837));
  inv1   g0522(.a(n837), .O(n838));
  nor2   g0523(.a(n838), .b(G1486), .O(n839));
  inv1   g0524(.a(G1486), .O(n840));
  nor2   g0525(.a(n837), .b(n840), .O(n841));
  nor2   g0526(.a(n841), .b(n839), .O(n842));
  inv1   g0527(.a(n842), .O(n843));
  nor2   g0528(.a(n843), .b(n835), .O(n844));
  inv1   g0529(.a(n844), .O(n845));
  nor2   g0530(.a(n845), .b(n797), .O(n846));
  inv1   g0531(.a(n809), .O(n847));
  nor2   g0532(.a(n847), .b(n805), .O(n848));
  nor2   g0533(.a(n848), .b(n801), .O(n849));
  inv1   g0534(.a(n849), .O(n850));
  nor2   g0535(.a(n850), .b(n827), .O(n851));
  nor2   g0536(.a(n851), .b(n829), .O(n852));
  nor2   g0537(.a(n852), .b(n819), .O(n853));
  nor2   g0538(.a(n853), .b(n821), .O(n854));
  inv1   g0539(.a(n854), .O(n855));
  nor2   g0540(.a(n855), .b(n841), .O(n856));
  nor2   g0541(.a(n856), .b(n839), .O(n857));
  inv1   g0542(.a(n857), .O(n858));
  nor2   g0543(.a(n858), .b(n846), .O(n859));
  nor2   g0544(.a(n859), .b(n393), .O(n860));
  nor2   g0545(.a(n860), .b(G38), .O(n861));
  inv1   g0546(.a(n859), .O(n862));
  inv1   g0547(.a(n387), .O(n863));
  nor2   g0548(.a(n863), .b(n388), .O(n864));
  inv1   g0549(.a(n864), .O(n865));
  nor2   g0550(.a(n865), .b(n862), .O(n866));
  nor2   g0551(.a(n866), .b(n861), .O(G246));
  inv1   g0552(.a(G38), .O(n868));
  nor2   g0553(.a(G2204), .b(G1455), .O(n869));
  inv1   g0554(.a(n869), .O(n870));
  nor2   g0555(.a(n870), .b(n386), .O(n871));
  nor2   g0556(.a(n871), .b(n868), .O(n872));
  inv1   g0557(.a(G206), .O(n873));
  nor2   g0558(.a(n873), .b(n397), .O(n874));
  nor2   g0559(.a(n874), .b(n518), .O(n875));
  nor2   g0560(.a(G3711), .b(n397), .O(n876));
  inv1   g0561(.a(G76), .O(n877));
  nor2   g0562(.a(n877), .b(G18), .O(n878));
  nor2   g0563(.a(n878), .b(n876), .O(n879));
  nor2   g0564(.a(n879), .b(n875), .O(n880));
  inv1   g0565(.a(G207), .O(n881));
  nor2   g0566(.a(n881), .b(n397), .O(n882));
  nor2   g0567(.a(n882), .b(n527), .O(n883));
  inv1   g0568(.a(n883), .O(n884));
  nor2   g0569(.a(G3705), .b(n397), .O(n885));
  inv1   g0570(.a(G74), .O(n886));
  nor2   g0571(.a(n886), .b(G18), .O(n887));
  nor2   g0572(.a(n887), .b(n885), .O(n888));
  inv1   g0573(.a(n888), .O(n889));
  nor2   g0574(.a(n889), .b(n884), .O(n890));
  nor2   g0575(.a(n888), .b(n883), .O(n891));
  inv1   g0576(.a(G70), .O(n892));
  nor2   g0577(.a(n892), .b(G18), .O(n893));
  nor2   g0578(.a(n893), .b(G89), .O(n894));
  inv1   g0579(.a(G89), .O(n895));
  nor2   g0580(.a(G70), .b(G18), .O(n896));
  nor2   g0581(.a(n896), .b(n895), .O(n897));
  nor2   g0582(.a(n897), .b(G41), .O(n898));
  nor2   g0583(.a(n898), .b(n894), .O(n899));
  nor2   g0584(.a(n899), .b(n891), .O(n900));
  nor2   g0585(.a(n900), .b(n890), .O(n901));
  nor2   g0586(.a(n901), .b(n880), .O(n902));
  inv1   g0587(.a(n875), .O(n903));
  inv1   g0588(.a(n879), .O(n904));
  nor2   g0589(.a(n904), .b(n903), .O(n905));
  inv1   g0590(.a(G205), .O(n906));
  nor2   g0591(.a(n906), .b(n397), .O(n907));
  nor2   g0592(.a(n907), .b(n504), .O(n908));
  inv1   g0593(.a(n908), .O(n909));
  nor2   g0594(.a(G3717), .b(n397), .O(n910));
  inv1   g0595(.a(G75), .O(n911));
  nor2   g0596(.a(n911), .b(G18), .O(n912));
  nor2   g0597(.a(n912), .b(n910), .O(n913));
  inv1   g0598(.a(n913), .O(n914));
  nor2   g0599(.a(n914), .b(n909), .O(n915));
  nor2   g0600(.a(n915), .b(n905), .O(n916));
  inv1   g0601(.a(n916), .O(n917));
  nor2   g0602(.a(n917), .b(n902), .O(n918));
  nor2   g0603(.a(n913), .b(n908), .O(n919));
  inv1   g0604(.a(G204), .O(n920));
  nor2   g0605(.a(n920), .b(n397), .O(n921));
  nor2   g0606(.a(n921), .b(n493), .O(n922));
  nor2   g0607(.a(G3723), .b(n397), .O(n923));
  inv1   g0608(.a(G73), .O(n924));
  nor2   g0609(.a(n924), .b(G18), .O(n925));
  nor2   g0610(.a(n925), .b(n923), .O(n926));
  nor2   g0611(.a(n926), .b(n922), .O(n927));
  nor2   g0612(.a(n927), .b(n919), .O(n928));
  inv1   g0613(.a(n928), .O(n929));
  nor2   g0614(.a(n929), .b(n918), .O(n930));
  inv1   g0615(.a(G200), .O(n931));
  nor2   g0616(.a(n931), .b(n397), .O(n932));
  nor2   g0617(.a(n932), .b(n467), .O(n933));
  nor2   g0618(.a(G3749), .b(n397), .O(n934));
  inv1   g0619(.a(G56), .O(n935));
  nor2   g0620(.a(n935), .b(G18), .O(n936));
  nor2   g0621(.a(n936), .b(n934), .O(n937));
  nor2   g0622(.a(n937), .b(n933), .O(n938));
  inv1   g0623(.a(G201), .O(n939));
  nor2   g0624(.a(n939), .b(n397), .O(n940));
  nor2   g0625(.a(n940), .b(n478), .O(n941));
  nor2   g0626(.a(G3743), .b(n397), .O(n942));
  inv1   g0627(.a(G55), .O(n943));
  nor2   g0628(.a(n943), .b(G18), .O(n944));
  nor2   g0629(.a(n944), .b(n942), .O(n945));
  nor2   g0630(.a(n945), .b(n941), .O(n946));
  nor2   g0631(.a(n946), .b(n938), .O(n947));
  inv1   g0632(.a(n947), .O(n948));
  inv1   g0633(.a(n933), .O(n949));
  inv1   g0634(.a(n937), .O(n950));
  nor2   g0635(.a(n950), .b(n949), .O(n951));
  inv1   g0636(.a(n941), .O(n952));
  inv1   g0637(.a(n945), .O(n953));
  nor2   g0638(.a(n953), .b(n952), .O(n954));
  nor2   g0639(.a(n954), .b(n951), .O(n955));
  inv1   g0640(.a(n955), .O(n956));
  nor2   g0641(.a(n956), .b(n948), .O(n957));
  inv1   g0642(.a(n957), .O(n958));
  inv1   g0643(.a(G203), .O(n959));
  nor2   g0644(.a(n959), .b(n397), .O(n960));
  nor2   g0645(.a(n960), .b(n443), .O(n961));
  nor2   g0646(.a(G3729), .b(n397), .O(n962));
  inv1   g0647(.a(G53), .O(n963));
  nor2   g0648(.a(n963), .b(G18), .O(n964));
  nor2   g0649(.a(n964), .b(n962), .O(n965));
  nor2   g0650(.a(n965), .b(n961), .O(n966));
  inv1   g0651(.a(G202), .O(n967));
  nor2   g0652(.a(n967), .b(n397), .O(n968));
  nor2   g0653(.a(n968), .b(n454), .O(n969));
  nor2   g0654(.a(G3737), .b(n397), .O(n970));
  inv1   g0655(.a(G54), .O(n971));
  nor2   g0656(.a(n971), .b(G18), .O(n972));
  nor2   g0657(.a(n972), .b(n970), .O(n973));
  nor2   g0658(.a(n973), .b(n969), .O(n974));
  nor2   g0659(.a(n974), .b(n966), .O(n975));
  inv1   g0660(.a(n975), .O(n976));
  inv1   g0661(.a(n961), .O(n977));
  inv1   g0662(.a(n965), .O(n978));
  nor2   g0663(.a(n978), .b(n977), .O(n979));
  inv1   g0664(.a(n922), .O(n980));
  inv1   g0665(.a(n926), .O(n981));
  nor2   g0666(.a(n981), .b(n980), .O(n982));
  inv1   g0667(.a(n969), .O(n983));
  inv1   g0668(.a(n973), .O(n984));
  nor2   g0669(.a(n984), .b(n983), .O(n985));
  nor2   g0670(.a(n985), .b(n982), .O(n986));
  inv1   g0671(.a(n986), .O(n987));
  nor2   g0672(.a(n987), .b(n979), .O(n988));
  inv1   g0673(.a(n988), .O(n989));
  nor2   g0674(.a(n989), .b(n976), .O(n990));
  inv1   g0675(.a(n990), .O(n991));
  nor2   g0676(.a(n991), .b(n958), .O(n992));
  inv1   g0677(.a(n992), .O(n993));
  nor2   g0678(.a(n993), .b(n930), .O(n994));
  nor2   g0679(.a(n951), .b(n947), .O(n995));
  nor2   g0680(.a(n985), .b(n975), .O(n996));
  inv1   g0681(.a(n996), .O(n997));
  nor2   g0682(.a(n997), .b(n958), .O(n998));
  nor2   g0683(.a(n998), .b(n995), .O(n999));
  inv1   g0684(.a(n999), .O(n1000));
  nor2   g0685(.a(n1000), .b(n994), .O(n1001));
  inv1   g0686(.a(G194), .O(n1002));
  nor2   g0687(.a(n1002), .b(n397), .O(n1003));
  nor2   g0688(.a(n1003), .b(n619), .O(n1004));
  nor2   g0689(.a(G4410), .b(n397), .O(n1005));
  inv1   g0690(.a(G81), .O(n1006));
  nor2   g0691(.a(n1006), .b(G18), .O(n1007));
  nor2   g0692(.a(n1007), .b(n1005), .O(n1008));
  nor2   g0693(.a(n1008), .b(n1004), .O(n1009));
  inv1   g0694(.a(G195), .O(n1010));
  nor2   g0695(.a(n1010), .b(n397), .O(n1011));
  nor2   g0696(.a(n1011), .b(n656), .O(n1012));
  nor2   g0697(.a(G4405), .b(n397), .O(n1013));
  inv1   g0698(.a(G59), .O(n1014));
  nor2   g0699(.a(n1014), .b(G18), .O(n1015));
  nor2   g0700(.a(n1015), .b(n1013), .O(n1016));
  nor2   g0701(.a(n1016), .b(n1012), .O(n1017));
  nor2   g0702(.a(n1017), .b(n1009), .O(n1018));
  inv1   g0703(.a(n1018), .O(n1019));
  inv1   g0704(.a(G196), .O(n1020));
  nor2   g0705(.a(n1020), .b(n397), .O(n1021));
  nor2   g0706(.a(n1021), .b(n632), .O(n1022));
  inv1   g0707(.a(n1022), .O(n1023));
  nor2   g0708(.a(G4400), .b(n397), .O(n1024));
  inv1   g0709(.a(G78), .O(n1025));
  nor2   g0710(.a(n1025), .b(G18), .O(n1026));
  nor2   g0711(.a(n1026), .b(n1024), .O(n1027));
  inv1   g0712(.a(n1027), .O(n1028));
  nor2   g0713(.a(n1028), .b(n1023), .O(n1029));
  inv1   g0714(.a(G193), .O(n1030));
  nor2   g0715(.a(n1030), .b(n397), .O(n1031));
  nor2   g0716(.a(n1031), .b(n608), .O(n1032));
  nor2   g0717(.a(G4415), .b(n397), .O(n1033));
  inv1   g0718(.a(G80), .O(n1034));
  nor2   g0719(.a(n1034), .b(G18), .O(n1035));
  nor2   g0720(.a(n1035), .b(n1033), .O(n1036));
  nor2   g0721(.a(n1036), .b(n1032), .O(n1037));
  nor2   g0722(.a(n1037), .b(n1029), .O(n1038));
  inv1   g0723(.a(n1038), .O(n1039));
  nor2   g0724(.a(n1039), .b(n1019), .O(n1040));
  inv1   g0725(.a(n1040), .O(n1041));
  inv1   g0726(.a(n1004), .O(n1042));
  inv1   g0727(.a(n1008), .O(n1043));
  nor2   g0728(.a(n1043), .b(n1042), .O(n1044));
  inv1   g0729(.a(n1012), .O(n1045));
  inv1   g0730(.a(n1016), .O(n1046));
  nor2   g0731(.a(n1046), .b(n1045), .O(n1047));
  nor2   g0732(.a(n1047), .b(n1044), .O(n1048));
  inv1   g0733(.a(n1048), .O(n1049));
  nor2   g0734(.a(n1027), .b(n1022), .O(n1050));
  inv1   g0735(.a(G187), .O(n1051));
  nor2   g0736(.a(n1051), .b(n397), .O(n1052));
  nor2   g0737(.a(n1052), .b(n643), .O(n1053));
  nor2   g0738(.a(G4394), .b(n397), .O(n1054));
  inv1   g0739(.a(G77), .O(n1055));
  nor2   g0740(.a(n1055), .b(G18), .O(n1056));
  nor2   g0741(.a(n1056), .b(n1054), .O(n1057));
  nor2   g0742(.a(n1057), .b(n1053), .O(n1058));
  nor2   g0743(.a(n1058), .b(n1050), .O(n1059));
  inv1   g0744(.a(n1059), .O(n1060));
  inv1   g0745(.a(n1032), .O(n1061));
  inv1   g0746(.a(n1036), .O(n1062));
  nor2   g0747(.a(n1062), .b(n1061), .O(n1063));
  inv1   g0748(.a(n1053), .O(n1064));
  inv1   g0749(.a(n1057), .O(n1065));
  nor2   g0750(.a(n1065), .b(n1064), .O(n1066));
  nor2   g0751(.a(n1066), .b(n1063), .O(n1067));
  inv1   g0752(.a(n1067), .O(n1068));
  nor2   g0753(.a(n1068), .b(n1060), .O(n1069));
  inv1   g0754(.a(n1069), .O(n1070));
  nor2   g0755(.a(n1070), .b(n1049), .O(n1071));
  inv1   g0756(.a(n1071), .O(n1072));
  nor2   g0757(.a(n1072), .b(n1041), .O(n1073));
  inv1   g0758(.a(n1073), .O(n1074));
  nor2   g0759(.a(n1074), .b(n1001), .O(n1075));
  nor2   g0760(.a(n1059), .b(n1029), .O(n1076));
  nor2   g0761(.a(n1076), .b(n1017), .O(n1077));
  nor2   g0762(.a(n1077), .b(n1049), .O(n1078));
  nor2   g0763(.a(n1037), .b(n1009), .O(n1079));
  inv1   g0764(.a(n1079), .O(n1080));
  nor2   g0765(.a(n1080), .b(n1078), .O(n1081));
  nor2   g0766(.a(n1081), .b(n1063), .O(n1082));
  nor2   g0767(.a(n1082), .b(n1075), .O(n1083));
  inv1   g0768(.a(G190), .O(n1084));
  nor2   g0769(.a(n1084), .b(n397), .O(n1085));
  nor2   g0770(.a(n1085), .b(n566), .O(n1086));
  inv1   g0771(.a(n1086), .O(n1087));
  nor2   g0772(.a(G4432), .b(n397), .O(n1088));
  inv1   g0773(.a(G61), .O(n1089));
  nor2   g0774(.a(n1089), .b(G18), .O(n1090));
  nor2   g0775(.a(n1090), .b(n1088), .O(n1091));
  inv1   g0776(.a(n1091), .O(n1092));
  nor2   g0777(.a(n1092), .b(n1087), .O(n1093));
  inv1   g0778(.a(G189), .O(n1094));
  nor2   g0779(.a(n1094), .b(n397), .O(n1095));
  nor2   g0780(.a(n1095), .b(n554), .O(n1096));
  nor2   g0781(.a(G4437), .b(n397), .O(n1097));
  inv1   g0782(.a(G62), .O(n1098));
  nor2   g0783(.a(n1098), .b(G18), .O(n1099));
  nor2   g0784(.a(n1099), .b(n1097), .O(n1100));
  nor2   g0785(.a(n1100), .b(n1096), .O(n1101));
  inv1   g0786(.a(n1096), .O(n1102));
  inv1   g0787(.a(n1100), .O(n1103));
  nor2   g0788(.a(n1103), .b(n1102), .O(n1104));
  nor2   g0789(.a(n1104), .b(n1101), .O(n1105));
  inv1   g0790(.a(n1105), .O(n1106));
  nor2   g0791(.a(n1106), .b(n1093), .O(n1107));
  inv1   g0792(.a(n1107), .O(n1108));
  nor2   g0793(.a(n1091), .b(n1086), .O(n1109));
  inv1   g0794(.a(G191), .O(n1110));
  nor2   g0795(.a(n1110), .b(n397), .O(n1111));
  nor2   g0796(.a(n1111), .b(n573), .O(n1112));
  nor2   g0797(.a(G4427), .b(n397), .O(n1113));
  inv1   g0798(.a(G60), .O(n1114));
  nor2   g0799(.a(n1114), .b(G18), .O(n1115));
  nor2   g0800(.a(n1115), .b(n1113), .O(n1116));
  nor2   g0801(.a(n1116), .b(n1112), .O(n1117));
  nor2   g0802(.a(n1117), .b(n1109), .O(n1118));
  inv1   g0803(.a(n1118), .O(n1119));
  inv1   g0804(.a(n1112), .O(n1120));
  inv1   g0805(.a(n1116), .O(n1121));
  nor2   g0806(.a(n1121), .b(n1120), .O(n1122));
  nor2   g0807(.a(n1122), .b(n1119), .O(n1123));
  inv1   g0808(.a(n1123), .O(n1124));
  nor2   g0809(.a(n1124), .b(n1108), .O(n1125));
  inv1   g0810(.a(n1125), .O(n1126));
  inv1   g0811(.a(G192), .O(n1127));
  nor2   g0812(.a(n1127), .b(n397), .O(n1128));
  nor2   g0813(.a(n1128), .b(n584), .O(n1129));
  inv1   g0814(.a(n1129), .O(n1130));
  nor2   g0815(.a(G4420), .b(n397), .O(n1131));
  inv1   g0816(.a(G79), .O(n1132));
  nor2   g0817(.a(n1132), .b(G18), .O(n1133));
  nor2   g0818(.a(n1133), .b(n1131), .O(n1134));
  inv1   g0819(.a(n1134), .O(n1135));
  nor2   g0820(.a(n1135), .b(n1130), .O(n1136));
  nor2   g0821(.a(n1134), .b(n1129), .O(n1137));
  nor2   g0822(.a(n1137), .b(n1136), .O(n1138));
  inv1   g0823(.a(n1138), .O(n1139));
  nor2   g0824(.a(n1139), .b(n1126), .O(n1140));
  inv1   g0825(.a(n1140), .O(n1141));
  nor2   g0826(.a(n1141), .b(n1083), .O(n1142));
  inv1   g0827(.a(n1137), .O(n1143));
  nor2   g0828(.a(n1143), .b(n1126), .O(n1144));
  nor2   g0829(.a(n1118), .b(n1108), .O(n1145));
  nor2   g0830(.a(n1145), .b(n1101), .O(n1146));
  inv1   g0831(.a(n1146), .O(n1147));
  nor2   g0832(.a(n1147), .b(n1144), .O(n1148));
  inv1   g0833(.a(n1148), .O(n1149));
  nor2   g0834(.a(n1149), .b(n1142), .O(n1150));
  nor2   g0835(.a(G173), .b(n397), .O(n1151));
  nor2   g0836(.a(n1151), .b(n396), .O(n1152));
  inv1   g0837(.a(G110), .O(n1153));
  nor2   g0838(.a(n1153), .b(G18), .O(n1154));
  nor2   g0839(.a(G2256), .b(n397), .O(n1155));
  nor2   g0840(.a(n1155), .b(n1154), .O(n1156));
  inv1   g0841(.a(n1156), .O(n1157));
  nor2   g0842(.a(n1157), .b(n1152), .O(n1158));
  nor2   g0843(.a(G174), .b(n397), .O(n1159));
  nor2   g0844(.a(n1159), .b(n396), .O(n1160));
  inv1   g0845(.a(G109), .O(n1161));
  nor2   g0846(.a(n1161), .b(G18), .O(n1162));
  nor2   g0847(.a(G2253), .b(n397), .O(n1163));
  nor2   g0848(.a(n1163), .b(n1162), .O(n1164));
  inv1   g0849(.a(n1164), .O(n1165));
  nor2   g0850(.a(n1165), .b(n1160), .O(n1166));
  nor2   g0851(.a(n1166), .b(n1158), .O(n1167));
  inv1   g0852(.a(n1167), .O(n1168));
  nor2   g0853(.a(G175), .b(n397), .O(n1169));
  nor2   g0854(.a(n1169), .b(n396), .O(n1170));
  inv1   g0855(.a(n1170), .O(n1171));
  inv1   g0856(.a(G86), .O(n1172));
  nor2   g0857(.a(n1172), .b(G18), .O(n1173));
  nor2   g0858(.a(G2247), .b(n397), .O(n1174));
  nor2   g0859(.a(n1174), .b(n1173), .O(n1175));
  nor2   g0860(.a(n1175), .b(n1171), .O(n1176));
  inv1   g0861(.a(n1160), .O(n1177));
  nor2   g0862(.a(n1164), .b(n1177), .O(n1178));
  nor2   g0863(.a(n1178), .b(n1176), .O(n1179));
  inv1   g0864(.a(n1179), .O(n1180));
  nor2   g0865(.a(n1180), .b(n1168), .O(n1181));
  inv1   g0866(.a(n1181), .O(n1182));
  nor2   g0867(.a(G177), .b(n397), .O(n1183));
  nor2   g0868(.a(n1183), .b(n396), .O(n1184));
  inv1   g0869(.a(n1184), .O(n1185));
  inv1   g0870(.a(G64), .O(n1186));
  nor2   g0871(.a(n1186), .b(G18), .O(n1187));
  nor2   g0872(.a(G2236), .b(n397), .O(n1188));
  nor2   g0873(.a(n1188), .b(n1187), .O(n1189));
  nor2   g0874(.a(n1189), .b(n1185), .O(n1190));
  inv1   g0875(.a(G178), .O(n1191));
  nor2   g0876(.a(n1191), .b(n397), .O(n1192));
  nor2   g0877(.a(n1192), .b(n715), .O(n1193));
  inv1   g0878(.a(G85), .O(n1194));
  nor2   g0879(.a(n1194), .b(G18), .O(n1195));
  nor2   g0880(.a(G2230), .b(n397), .O(n1196));
  nor2   g0881(.a(n1196), .b(n1195), .O(n1197));
  nor2   g0882(.a(n1197), .b(n1193), .O(n1198));
  nor2   g0883(.a(n1198), .b(n1190), .O(n1199));
  inv1   g0884(.a(n1199), .O(n1200));
  inv1   g0885(.a(G171), .O(n1201));
  nor2   g0886(.a(n1201), .b(n397), .O(n1202));
  nor2   g0887(.a(n1202), .b(n750), .O(n1203));
  inv1   g0888(.a(G65), .O(n1204));
  nor2   g0889(.a(n1204), .b(G18), .O(n1205));
  nor2   g0890(.a(G2211), .b(n397), .O(n1206));
  nor2   g0891(.a(n1206), .b(n1205), .O(n1207));
  nor2   g0892(.a(n1207), .b(n1203), .O(n1208));
  inv1   g0893(.a(G180), .O(n1209));
  nor2   g0894(.a(n1209), .b(n397), .O(n1210));
  nor2   g0895(.a(n1210), .b(n739), .O(n1211));
  inv1   g0896(.a(G83), .O(n1212));
  nor2   g0897(.a(n1212), .b(G18), .O(n1213));
  nor2   g0898(.a(G2218), .b(n397), .O(n1214));
  nor2   g0899(.a(n1214), .b(n1213), .O(n1215));
  nor2   g0900(.a(n1215), .b(n1211), .O(n1216));
  nor2   g0901(.a(n1216), .b(n1208), .O(n1217));
  inv1   g0902(.a(n1217), .O(n1218));
  nor2   g0903(.a(n1218), .b(n1200), .O(n1219));
  inv1   g0904(.a(n1219), .O(n1220));
  nor2   g0905(.a(n1220), .b(n1182), .O(n1221));
  inv1   g0906(.a(n1221), .O(n1222));
  inv1   g0907(.a(G179), .O(n1223));
  nor2   g0908(.a(n1223), .b(n397), .O(n1224));
  nor2   g0909(.a(n1224), .b(n726), .O(n1225));
  inv1   g0910(.a(n1225), .O(n1226));
  inv1   g0911(.a(G84), .O(n1227));
  nor2   g0912(.a(n1227), .b(G18), .O(n1228));
  nor2   g0913(.a(G2224), .b(n397), .O(n1229));
  nor2   g0914(.a(n1229), .b(n1228), .O(n1230));
  inv1   g0915(.a(n1230), .O(n1231));
  nor2   g0916(.a(n1231), .b(n1226), .O(n1232));
  nor2   g0917(.a(n1230), .b(n1225), .O(n1233));
  inv1   g0918(.a(n1211), .O(n1234));
  inv1   g0919(.a(n1215), .O(n1235));
  nor2   g0920(.a(n1235), .b(n1234), .O(n1236));
  nor2   g0921(.a(n1236), .b(n1233), .O(n1237));
  inv1   g0922(.a(n1237), .O(n1238));
  nor2   g0923(.a(n1238), .b(n1232), .O(n1239));
  inv1   g0924(.a(n1239), .O(n1240));
  inv1   g0925(.a(n1189), .O(n1241));
  nor2   g0926(.a(n1241), .b(n1184), .O(n1242));
  nor2   g0927(.a(G176), .b(n397), .O(n1243));
  nor2   g0928(.a(n1243), .b(n396), .O(n1244));
  inv1   g0929(.a(n1244), .O(n1245));
  inv1   g0930(.a(G63), .O(n1246));
  nor2   g0931(.a(n1246), .b(G18), .O(n1247));
  nor2   g0932(.a(G2239), .b(n397), .O(n1248));
  nor2   g0933(.a(n1248), .b(n1247), .O(n1249));
  nor2   g0934(.a(n1249), .b(n1245), .O(n1250));
  inv1   g0935(.a(n1249), .O(n1251));
  nor2   g0936(.a(n1251), .b(n1244), .O(n1252));
  nor2   g0937(.a(n1252), .b(n1250), .O(n1253));
  inv1   g0938(.a(n1253), .O(n1254));
  nor2   g0939(.a(n1254), .b(n1242), .O(n1255));
  inv1   g0940(.a(n1255), .O(n1256));
  inv1   g0941(.a(n1152), .O(n1257));
  nor2   g0942(.a(n1156), .b(n1257), .O(n1258));
  inv1   g0943(.a(n1175), .O(n1259));
  nor2   g0944(.a(n1259), .b(n1170), .O(n1260));
  nor2   g0945(.a(n1260), .b(n1258), .O(n1261));
  inv1   g0946(.a(n1261), .O(n1262));
  inv1   g0947(.a(n1193), .O(n1263));
  inv1   g0948(.a(n1197), .O(n1264));
  nor2   g0949(.a(n1264), .b(n1263), .O(n1265));
  inv1   g0950(.a(n1203), .O(n1266));
  inv1   g0951(.a(n1207), .O(n1267));
  nor2   g0952(.a(n1267), .b(n1266), .O(n1268));
  nor2   g0953(.a(n1268), .b(n1265), .O(n1269));
  inv1   g0954(.a(n1269), .O(n1270));
  nor2   g0955(.a(n1270), .b(n1262), .O(n1271));
  inv1   g0956(.a(n1271), .O(n1272));
  nor2   g0957(.a(n1272), .b(n1256), .O(n1273));
  inv1   g0958(.a(n1273), .O(n1274));
  nor2   g0959(.a(n1274), .b(n1240), .O(n1275));
  inv1   g0960(.a(n1275), .O(n1276));
  nor2   g0961(.a(n1276), .b(n1222), .O(n1277));
  inv1   g0962(.a(n1277), .O(n1278));
  nor2   g0963(.a(n1278), .b(n1150), .O(n1279));
  nor2   g0964(.a(n1265), .b(n1198), .O(n1280));
  inv1   g0965(.a(n1280), .O(n1281));
  nor2   g0966(.a(n1281), .b(n1217), .O(n1282));
  inv1   g0967(.a(n1282), .O(n1283));
  nor2   g0968(.a(n1283), .b(n1240), .O(n1284));
  inv1   g0969(.a(n1233), .O(n1285));
  nor2   g0970(.a(n1281), .b(n1285), .O(n1286));
  nor2   g0971(.a(n1286), .b(n1200), .O(n1287));
  inv1   g0972(.a(n1287), .O(n1288));
  nor2   g0973(.a(n1288), .b(n1284), .O(n1289));
  nor2   g0974(.a(n1289), .b(n1256), .O(n1290));
  nor2   g0975(.a(n1290), .b(n1250), .O(n1291));
  nor2   g0976(.a(n1291), .b(n1260), .O(n1292));
  nor2   g0977(.a(n1292), .b(n1180), .O(n1293));
  nor2   g0978(.a(n1293), .b(n1168), .O(n1294));
  nor2   g0979(.a(n1294), .b(n1258), .O(n1295));
  inv1   g0980(.a(n1295), .O(n1296));
  nor2   g0981(.a(n1296), .b(n1279), .O(n1297));
  nor2   g0982(.a(G167), .b(n397), .O(n1298));
  nor2   g0983(.a(n1298), .b(n396), .O(n1299));
  inv1   g0984(.a(n1299), .O(n1300));
  inv1   g0985(.a(G112), .O(n1301));
  nor2   g0986(.a(n1301), .b(G18), .O(n1302));
  nor2   g0987(.a(G1480), .b(n397), .O(n1303));
  nor2   g0988(.a(n1303), .b(n1302), .O(n1304));
  nor2   g0989(.a(n1304), .b(n1300), .O(n1305));
  nor2   g0990(.a(G168), .b(n397), .O(n1306));
  nor2   g0991(.a(n1306), .b(n396), .O(n1307));
  inv1   g0992(.a(G87), .O(n1308));
  nor2   g0993(.a(n1308), .b(G18), .O(n1309));
  nor2   g0994(.a(G106), .b(n397), .O(n1310));
  nor2   g0995(.a(n1310), .b(n1309), .O(n1311));
  inv1   g0996(.a(n1311), .O(n1312));
  nor2   g0997(.a(n1312), .b(n1307), .O(n1313));
  nor2   g0998(.a(n1313), .b(n1305), .O(n1314));
  inv1   g0999(.a(n1314), .O(n1315));
  inv1   g1000(.a(n1304), .O(n1316));
  nor2   g1001(.a(n1316), .b(n1299), .O(n1317));
  inv1   g1002(.a(n1307), .O(n1318));
  nor2   g1003(.a(n1311), .b(n1318), .O(n1319));
  nor2   g1004(.a(n1319), .b(n1317), .O(n1320));
  inv1   g1005(.a(n1320), .O(n1321));
  nor2   g1006(.a(n1321), .b(n1315), .O(n1322));
  inv1   g1007(.a(n1322), .O(n1323));
  nor2   g1008(.a(G169), .b(n397), .O(n1324));
  nor2   g1009(.a(n1324), .b(n396), .O(n1325));
  inv1   g1010(.a(G111), .O(n1326));
  nor2   g1011(.a(n1326), .b(G18), .O(n1327));
  nor2   g1012(.a(G1469), .b(n397), .O(n1328));
  nor2   g1013(.a(n1328), .b(n1327), .O(n1329));
  inv1   g1014(.a(n1329), .O(n1330));
  nor2   g1015(.a(n1330), .b(n1325), .O(n1331));
  inv1   g1016(.a(n1325), .O(n1332));
  nor2   g1017(.a(n1329), .b(n1332), .O(n1333));
  nor2   g1018(.a(n1333), .b(n1331), .O(n1334));
  inv1   g1019(.a(n1334), .O(n1335));
  nor2   g1020(.a(n1335), .b(n1323), .O(n1336));
  inv1   g1021(.a(n1336), .O(n1337));
  nor2   g1022(.a(G166), .b(n397), .O(n1338));
  nor2   g1023(.a(n1338), .b(n396), .O(n1339));
  inv1   g1024(.a(n1339), .O(n1340));
  inv1   g1025(.a(G88), .O(n1341));
  nor2   g1026(.a(n1341), .b(G18), .O(n1342));
  nor2   g1027(.a(G1486), .b(n397), .O(n1343));
  nor2   g1028(.a(n1343), .b(n1342), .O(n1344));
  nor2   g1029(.a(n1344), .b(n1340), .O(n1345));
  inv1   g1030(.a(G113), .O(n1346));
  nor2   g1031(.a(n1346), .b(G18), .O(n1347));
  nor2   g1032(.a(G1462), .b(n397), .O(n1348));
  nor2   g1033(.a(n1348), .b(n1347), .O(n1349));
  nor2   g1034(.a(n1349), .b(n396), .O(n1350));
  nor2   g1035(.a(n1350), .b(n1345), .O(n1351));
  inv1   g1036(.a(n1351), .O(n1352));
  inv1   g1037(.a(n1344), .O(n1353));
  nor2   g1038(.a(n1353), .b(n1339), .O(n1354));
  inv1   g1039(.a(n396), .O(n1355));
  inv1   g1040(.a(n1349), .O(n1356));
  nor2   g1041(.a(n1356), .b(n1355), .O(n1357));
  nor2   g1042(.a(n1357), .b(n1354), .O(n1358));
  inv1   g1043(.a(n1358), .O(n1359));
  nor2   g1044(.a(n1359), .b(n1352), .O(n1360));
  inv1   g1045(.a(n1360), .O(n1361));
  nor2   g1046(.a(n1361), .b(n1337), .O(n1362));
  inv1   g1047(.a(n1362), .O(n1363));
  nor2   g1048(.a(n1363), .b(n1297), .O(n1364));
  inv1   g1049(.a(n1350), .O(n1365));
  nor2   g1050(.a(n1365), .b(n1337), .O(n1366));
  inv1   g1051(.a(n1333), .O(n1367));
  nor2   g1052(.a(n1367), .b(n1323), .O(n1368));
  inv1   g1053(.a(n1319), .O(n1369));
  nor2   g1054(.a(n1369), .b(n1317), .O(n1370));
  nor2   g1055(.a(n1345), .b(n1305), .O(n1371));
  inv1   g1056(.a(n1371), .O(n1372));
  nor2   g1057(.a(n1372), .b(n1370), .O(n1373));
  inv1   g1058(.a(n1373), .O(n1374));
  nor2   g1059(.a(n1374), .b(n1368), .O(n1375));
  inv1   g1060(.a(n1375), .O(n1376));
  nor2   g1061(.a(n1376), .b(n1366), .O(n1377));
  nor2   g1062(.a(n1377), .b(n1354), .O(n1378));
  nor2   g1063(.a(n1378), .b(n1364), .O(n1379));
  inv1   g1064(.a(G1455), .O(n1380));
  inv1   g1065(.a(G2204), .O(n1381));
  nor2   g1066(.a(n1381), .b(n1380), .O(n1382));
  nor2   g1067(.a(n386), .b(G38), .O(n1383));
  inv1   g1068(.a(n1383), .O(n1384));
  nor2   g1069(.a(n1384), .b(n1382), .O(n1385));
  nor2   g1070(.a(n1385), .b(n1379), .O(n1386));
  nor2   g1071(.a(n1386), .b(n872), .O(n1387));
  inv1   g1072(.a(n1387), .O(G258));
  nor2   g1073(.a(n697), .b(n535), .O(n1389));
  nor2   g1074(.a(n1389), .b(n511), .O(n1390));
  nor2   g1075(.a(n1390), .b(n506), .O(n1391));
  nor2   g1076(.a(n1391), .b(n500), .O(n1392));
  inv1   g1077(.a(n1391), .O(n1393));
  nor2   g1078(.a(n1393), .b(n499), .O(n1394));
  nor2   g1079(.a(n1394), .b(n1392), .O(G388));
  inv1   g1080(.a(n1389), .O(n1396));
  nor2   g1081(.a(n1396), .b(n510), .O(n1397));
  nor2   g1082(.a(n1397), .b(n1390), .O(G391));
  nor2   g1083(.a(n382), .b(n375), .O(n1399));
  nor2   g1084(.a(n1399), .b(n690), .O(n1400));
  nor2   g1085(.a(n1400), .b(n531), .O(n1401));
  nor2   g1086(.a(n1401), .b(n694), .O(n1402));
  inv1   g1087(.a(n1401), .O(n1403));
  nor2   g1088(.a(n1403), .b(n693), .O(n1404));
  nor2   g1089(.a(n1404), .b(n1402), .O(G394));
  inv1   g1090(.a(n1399), .O(n1406));
  nor2   g1091(.a(n1406), .b(n689), .O(n1407));
  nor2   g1092(.a(n1407), .b(n1400), .O(G397));
  inv1   g1093(.a(n546), .O(n1409));
  inv1   g1094(.a(n544), .O(n1410));
  inv1   g1095(.a(n540), .O(n1411));
  nor2   g1096(.a(n699), .b(n1411), .O(n1412));
  nor2   g1097(.a(n1412), .b(n463), .O(n1413));
  nor2   g1098(.a(n1413), .b(n1410), .O(n1414));
  nor2   g1099(.a(n1414), .b(n485), .O(n1415));
  nor2   g1100(.a(n1415), .b(n1409), .O(n1416));
  nor2   g1101(.a(n1416), .b(n474), .O(n1417));
  inv1   g1102(.a(n1416), .O(n1418));
  nor2   g1103(.a(n1418), .b(n473), .O(n1419));
  nor2   g1104(.a(n1419), .b(n1417), .O(G376));
  inv1   g1105(.a(n1414), .O(n1421));
  nor2   g1106(.a(n1421), .b(n484), .O(n1422));
  nor2   g1107(.a(n1422), .b(n1415), .O(G379));
  nor2   g1108(.a(n1412), .b(n450), .O(n1424));
  nor2   g1109(.a(n460), .b(n445), .O(n1425));
  nor2   g1110(.a(n1425), .b(n543), .O(n1426));
  nor2   g1111(.a(n1426), .b(n1424), .O(n1427));
  nor2   g1112(.a(n1427), .b(n1413), .O(G382));
  inv1   g1113(.a(n1412), .O(n1429));
  nor2   g1114(.a(n1429), .b(n449), .O(n1430));
  nor2   g1115(.a(n1430), .b(n1424), .O(G385));
  nor2   g1116(.a(n620), .b(n595), .O(n1432));
  nor2   g1117(.a(n623), .b(n585), .O(n1433));
  nor2   g1118(.a(n1433), .b(n1432), .O(n1434));
  inv1   g1119(.a(n1434), .O(n1435));
  nor2   g1120(.a(n633), .b(n568), .O(n1436));
  nor2   g1121(.a(n636), .b(n567), .O(n1437));
  nor2   g1122(.a(n1437), .b(n1436), .O(n1438));
  nor2   g1123(.a(n1438), .b(n558), .O(n1439));
  inv1   g1124(.a(n1438), .O(n1440));
  nor2   g1125(.a(n1440), .b(n555), .O(n1441));
  nor2   g1126(.a(n1441), .b(n1439), .O(n1442));
  inv1   g1127(.a(n1442), .O(n1443));
  nor2   g1128(.a(n1443), .b(n577), .O(n1444));
  nor2   g1129(.a(n1442), .b(n574), .O(n1445));
  nor2   g1130(.a(n1445), .b(n1444), .O(n1446));
  inv1   g1131(.a(G227), .O(n1447));
  nor2   g1132(.a(n1447), .b(n397), .O(n1448));
  inv1   g1133(.a(G115), .O(n1449));
  nor2   g1134(.a(n1449), .b(G18), .O(n1450));
  nor2   g1135(.a(n1450), .b(n1448), .O(n1451));
  nor2   g1136(.a(n1451), .b(n612), .O(n1452));
  inv1   g1137(.a(n1451), .O(n1453));
  nor2   g1138(.a(n1453), .b(n609), .O(n1454));
  nor2   g1139(.a(n1454), .b(n1452), .O(n1455));
  inv1   g1140(.a(n1455), .O(n1456));
  nor2   g1141(.a(n1456), .b(n647), .O(n1457));
  nor2   g1142(.a(n1455), .b(n644), .O(n1458));
  nor2   g1143(.a(n1458), .b(n1457), .O(n1459));
  nor2   g1144(.a(n1459), .b(n660), .O(n1460));
  inv1   g1145(.a(n1459), .O(n1461));
  nor2   g1146(.a(n1461), .b(n657), .O(n1462));
  nor2   g1147(.a(n1462), .b(n1460), .O(n1463));
  inv1   g1148(.a(n1463), .O(n1464));
  nor2   g1149(.a(n1464), .b(n1446), .O(n1465));
  inv1   g1150(.a(n1446), .O(n1466));
  nor2   g1151(.a(n1463), .b(n1466), .O(n1467));
  nor2   g1152(.a(n1467), .b(n1465), .O(n1468));
  nor2   g1153(.a(n1468), .b(n1435), .O(n1469));
  inv1   g1154(.a(n1468), .O(n1470));
  nor2   g1155(.a(n1470), .b(n1434), .O(n1471));
  nor2   g1156(.a(n1471), .b(n1469), .O(n1472));
  nor2   g1157(.a(n528), .b(n497), .O(n1473));
  nor2   g1158(.a(n529), .b(n494), .O(n1474));
  nor2   g1159(.a(n1474), .b(n1473), .O(n1475));
  nor2   g1160(.a(n1475), .b(n482), .O(n1476));
  inv1   g1161(.a(n1475), .O(n1477));
  nor2   g1162(.a(n1477), .b(n479), .O(n1478));
  nor2   g1163(.a(n1478), .b(n1476), .O(n1479));
  inv1   g1164(.a(G239), .O(n1480));
  nor2   g1165(.a(n1480), .b(n397), .O(n1481));
  inv1   g1166(.a(G44), .O(n1482));
  nor2   g1167(.a(n1482), .b(G18), .O(n1483));
  nor2   g1168(.a(n1483), .b(n1481), .O(n1484));
  inv1   g1169(.a(n1484), .O(n1485));
  inv1   g1170(.a(G229), .O(n1486));
  nor2   g1171(.a(n1486), .b(n397), .O(n1487));
  nor2   g1172(.a(n1487), .b(n373), .O(n1488));
  nor2   g1173(.a(n1488), .b(n520), .O(n1489));
  inv1   g1174(.a(n1488), .O(n1490));
  nor2   g1175(.a(n1490), .b(n519), .O(n1491));
  nor2   g1176(.a(n1491), .b(n1489), .O(n1492));
  inv1   g1177(.a(n1492), .O(n1493));
  nor2   g1178(.a(n1493), .b(n1485), .O(n1494));
  nor2   g1179(.a(n1492), .b(n1484), .O(n1495));
  nor2   g1180(.a(n1495), .b(n1494), .O(n1496));
  nor2   g1181(.a(n505), .b(n471), .O(n1497));
  nor2   g1182(.a(n508), .b(n468), .O(n1498));
  nor2   g1183(.a(n1498), .b(n1497), .O(n1499));
  inv1   g1184(.a(n1499), .O(n1500));
  nor2   g1185(.a(n1500), .b(n458), .O(n1501));
  nor2   g1186(.a(n1499), .b(n455), .O(n1502));
  nor2   g1187(.a(n1502), .b(n1501), .O(n1503));
  nor2   g1188(.a(n1503), .b(n447), .O(n1504));
  inv1   g1189(.a(n1503), .O(n1505));
  nor2   g1190(.a(n1505), .b(n444), .O(n1506));
  nor2   g1191(.a(n1506), .b(n1504), .O(n1507));
  inv1   g1192(.a(n1507), .O(n1508));
  nor2   g1193(.a(n1508), .b(n1496), .O(n1509));
  inv1   g1194(.a(n1496), .O(n1510));
  nor2   g1195(.a(n1507), .b(n1510), .O(n1511));
  nor2   g1196(.a(n1511), .b(n1509), .O(n1512));
  nor2   g1197(.a(n1512), .b(n1479), .O(n1513));
  inv1   g1198(.a(n836), .O(n1514));
  nor2   g1199(.a(n1514), .b(n818), .O(n1515));
  inv1   g1200(.a(n816), .O(n1516));
  nor2   g1201(.a(n838), .b(n1516), .O(n1517));
  nor2   g1202(.a(n1517), .b(n1515), .O(n1518));
  inv1   g1203(.a(n1518), .O(n1519));
  nor2   g1204(.a(n396), .b(n397), .O(n1520));
  inv1   g1205(.a(n1520), .O(n1521));
  inv1   g1206(.a(G211), .O(n1522));
  inv1   g1207(.a(G212), .O(n1523));
  nor2   g1208(.a(n1523), .b(n1522), .O(n1524));
  nor2   g1209(.a(G212), .b(G211), .O(n1525));
  nor2   g1210(.a(n1525), .b(n1524), .O(n1526));
  inv1   g1211(.a(n1526), .O(n1527));
  nor2   g1212(.a(n1527), .b(n1521), .O(n1528));
  inv1   g1213(.a(n1528), .O(n1529));
  inv1   g1214(.a(n806), .O(n1530));
  inv1   g1215(.a(n798), .O(n1531));
  nor2   g1216(.a(n824), .b(n1531), .O(n1532));
  inv1   g1217(.a(n824), .O(n1533));
  nor2   g1218(.a(n1533), .b(n798), .O(n1534));
  nor2   g1219(.a(n1534), .b(n1532), .O(n1535));
  inv1   g1220(.a(n1535), .O(n1536));
  nor2   g1221(.a(n1536), .b(n1530), .O(n1537));
  nor2   g1222(.a(n1535), .b(n806), .O(n1538));
  nor2   g1223(.a(n1538), .b(n1537), .O(n1539));
  nor2   g1224(.a(n1539), .b(n1529), .O(n1540));
  nor2   g1225(.a(n1539), .b(n396), .O(n1541));
  nor2   g1226(.a(n1541), .b(n1528), .O(n1542));
  nor2   g1227(.a(n1542), .b(n1540), .O(n1543));
  nor2   g1228(.a(n1543), .b(n1519), .O(n1544));
  inv1   g1229(.a(n1543), .O(n1545));
  nor2   g1230(.a(n1545), .b(n1518), .O(n1546));
  nor2   g1231(.a(n1546), .b(n1544), .O(n1547));
  inv1   g1232(.a(n1479), .O(n1548));
  inv1   g1233(.a(n1512), .O(n1549));
  nor2   g1234(.a(n1549), .b(n1548), .O(n1550));
  nor2   g1235(.a(n1550), .b(n1547), .O(n1551));
  inv1   g1236(.a(n1551), .O(n1552));
  nor2   g1237(.a(n1552), .b(n1513), .O(n1553));
  inv1   g1238(.a(n1553), .O(n1554));
  nor2   g1239(.a(n1554), .b(n1472), .O(n1555));
  inv1   g1240(.a(n1555), .O(n1556));
  inv1   g1241(.a(G141), .O(n1557));
  nor2   g1242(.a(n1557), .b(G18), .O(n1558));
  inv1   g1243(.a(G161), .O(n1559));
  nor2   g1244(.a(n1559), .b(n397), .O(n1560));
  nor2   g1245(.a(n1560), .b(n1558), .O(n1561));
  nor2   g1246(.a(n1561), .b(n756), .O(n1562));
  inv1   g1247(.a(n1561), .O(n1563));
  nor2   g1248(.a(n1563), .b(n753), .O(n1564));
  nor2   g1249(.a(n1564), .b(n1562), .O(n1565));
  inv1   g1250(.a(n1565), .O(n1566));
  inv1   g1251(.a(n398), .O(n1567));
  nor2   g1252(.a(n428), .b(n1567), .O(n1568));
  inv1   g1253(.a(n407), .O(n1569));
  nor2   g1254(.a(n1569), .b(n400), .O(n1570));
  nor2   g1255(.a(n1570), .b(n1568), .O(n1571));
  nor2   g1256(.a(n1571), .b(n721), .O(n1572));
  inv1   g1257(.a(n1571), .O(n1573));
  nor2   g1258(.a(n1573), .b(n718), .O(n1574));
  nor2   g1259(.a(n1574), .b(n1572), .O(n1575));
  inv1   g1260(.a(n1575), .O(n1576));
  inv1   g1261(.a(n410), .O(n1577));
  nor2   g1262(.a(n420), .b(n1577), .O(n1578));
  inv1   g1263(.a(n418), .O(n1579));
  nor2   g1264(.a(n1579), .b(n412), .O(n1580));
  nor2   g1265(.a(n1580), .b(n1578), .O(n1581));
  nor2   g1266(.a(n1581), .b(n745), .O(n1582));
  inv1   g1267(.a(n1581), .O(n1583));
  nor2   g1268(.a(n1583), .b(n742), .O(n1584));
  nor2   g1269(.a(n1584), .b(n1582), .O(n1585));
  nor2   g1270(.a(n1585), .b(n732), .O(n1586));
  inv1   g1271(.a(n1585), .O(n1587));
  nor2   g1272(.a(n1587), .b(n729), .O(n1588));
  nor2   g1273(.a(n1588), .b(n1586), .O(n1589));
  inv1   g1274(.a(n1589), .O(n1590));
  nor2   g1275(.a(n1590), .b(n1576), .O(n1591));
  nor2   g1276(.a(n1589), .b(n1575), .O(n1592));
  nor2   g1277(.a(n1592), .b(n1591), .O(n1593));
  nor2   g1278(.a(n1593), .b(n766), .O(n1594));
  inv1   g1279(.a(n1593), .O(n1595));
  nor2   g1280(.a(n1595), .b(n765), .O(n1596));
  nor2   g1281(.a(n1596), .b(n1594), .O(n1597));
  inv1   g1282(.a(n1597), .O(n1598));
  nor2   g1283(.a(n1598), .b(n1566), .O(n1599));
  nor2   g1284(.a(n1597), .b(n1565), .O(n1600));
  nor2   g1285(.a(n1600), .b(n1599), .O(n1601));
  inv1   g1286(.a(n1601), .O(n1602));
  nor2   g1287(.a(n1602), .b(n1556), .O(n1603));
  inv1   g1288(.a(n1603), .O(G412));
  nor2   g1289(.a(n1197), .b(n1165), .O(n1605));
  nor2   g1290(.a(n1264), .b(n1164), .O(n1606));
  nor2   g1291(.a(n1606), .b(n1605), .O(n1607));
  inv1   g1292(.a(n1607), .O(n1608));
  nor2   g1293(.a(n1215), .b(n1157), .O(n1609));
  nor2   g1294(.a(n1235), .b(n1156), .O(n1610));
  nor2   g1295(.a(n1610), .b(n1609), .O(n1611));
  nor2   g1296(.a(n1611), .b(n1259), .O(n1612));
  inv1   g1297(.a(n1611), .O(n1613));
  nor2   g1298(.a(n1613), .b(n1175), .O(n1614));
  nor2   g1299(.a(n1614), .b(n1612), .O(n1615));
  inv1   g1300(.a(n1615), .O(n1616));
  nor2   g1301(.a(n1616), .b(n1251), .O(n1617));
  nor2   g1302(.a(n1615), .b(n1249), .O(n1618));
  nor2   g1303(.a(n1618), .b(n1617), .O(n1619));
  nor2   g1304(.a(n1619), .b(n1231), .O(n1620));
  inv1   g1305(.a(n1619), .O(n1621));
  nor2   g1306(.a(n1621), .b(n1230), .O(n1622));
  nor2   g1307(.a(n1622), .b(n1620), .O(n1623));
  inv1   g1308(.a(n1623), .O(n1624));
  nor2   g1309(.a(n1624), .b(n1608), .O(n1625));
  nor2   g1310(.a(n1623), .b(n1607), .O(n1626));
  nor2   g1311(.a(n1626), .b(n1625), .O(n1627));
  inv1   g1312(.a(n1627), .O(n1628));
  nor2   g1313(.a(G82), .b(G18), .O(n1629));
  inv1   g1314(.a(G2208), .O(n1630));
  nor2   g1315(.a(n1630), .b(n397), .O(n1631));
  nor2   g1316(.a(n1631), .b(n1629), .O(n1632));
  nor2   g1317(.a(n1632), .b(n1241), .O(n1633));
  inv1   g1318(.a(n1632), .O(n1634));
  nor2   g1319(.a(n1634), .b(n1189), .O(n1635));
  nor2   g1320(.a(n1635), .b(n1633), .O(n1636));
  nor2   g1321(.a(n1636), .b(n1207), .O(n1637));
  inv1   g1322(.a(n1636), .O(n1638));
  nor2   g1323(.a(n1638), .b(n1267), .O(n1639));
  nor2   g1324(.a(n1639), .b(n1637), .O(n1640));
  nor2   g1325(.a(n1640), .b(n1628), .O(n1641));
  inv1   g1326(.a(n1640), .O(n1642));
  nor2   g1327(.a(n1642), .b(n1627), .O(n1643));
  nor2   g1328(.a(n1643), .b(n1641), .O(n1644));
  nor2   g1329(.a(G4393), .b(n397), .O(n1645));
  inv1   g1330(.a(G58), .O(n1646));
  nor2   g1331(.a(n1646), .b(G18), .O(n1647));
  nor2   g1332(.a(n1647), .b(n1645), .O(n1648));
  nor2   g1333(.a(n1648), .b(n1135), .O(n1649));
  inv1   g1334(.a(n1648), .O(n1650));
  nor2   g1335(.a(n1650), .b(n1134), .O(n1651));
  nor2   g1336(.a(n1651), .b(n1649), .O(n1652));
  nor2   g1337(.a(n1652), .b(n1092), .O(n1653));
  inv1   g1338(.a(n1652), .O(n1654));
  nor2   g1339(.a(n1654), .b(n1091), .O(n1655));
  nor2   g1340(.a(n1655), .b(n1653), .O(n1656));
  nor2   g1341(.a(n1036), .b(n1043), .O(n1657));
  nor2   g1342(.a(n1062), .b(n1008), .O(n1658));
  nor2   g1343(.a(n1658), .b(n1657), .O(n1659));
  inv1   g1344(.a(n1659), .O(n1660));
  nor2   g1345(.a(n1660), .b(n1065), .O(n1661));
  nor2   g1346(.a(n1659), .b(n1057), .O(n1662));
  nor2   g1347(.a(n1662), .b(n1661), .O(n1663));
  nor2   g1348(.a(n1663), .b(n1046), .O(n1664));
  inv1   g1349(.a(n1663), .O(n1665));
  nor2   g1350(.a(n1665), .b(n1016), .O(n1666));
  nor2   g1351(.a(n1666), .b(n1664), .O(n1667));
  inv1   g1352(.a(n1667), .O(n1668));
  nor2   g1353(.a(n1668), .b(n1028), .O(n1669));
  nor2   g1354(.a(n1667), .b(n1027), .O(n1670));
  nor2   g1355(.a(n1670), .b(n1669), .O(n1671));
  inv1   g1356(.a(n1671), .O(n1672));
  nor2   g1357(.a(n1116), .b(n1103), .O(n1673));
  nor2   g1358(.a(n1121), .b(n1100), .O(n1674));
  nor2   g1359(.a(n1674), .b(n1673), .O(n1675));
  nor2   g1360(.a(n1675), .b(n1672), .O(n1676));
  inv1   g1361(.a(n1675), .O(n1677));
  nor2   g1362(.a(n1677), .b(n1671), .O(n1678));
  nor2   g1363(.a(n1678), .b(n1676), .O(n1679));
  nor2   g1364(.a(n1679), .b(n1656), .O(n1680));
  inv1   g1365(.a(n1656), .O(n1681));
  inv1   g1366(.a(n1679), .O(n1682));
  nor2   g1367(.a(n1682), .b(n1681), .O(n1683));
  nor2   g1368(.a(G1455), .b(G18), .O(n1684));
  nor2   g1369(.a(n388), .b(n397), .O(n1685));
  nor2   g1370(.a(n1685), .b(n1684), .O(n1686));
  nor2   g1371(.a(n1686), .b(n1316), .O(n1687));
  inv1   g1372(.a(n1686), .O(n1688));
  nor2   g1373(.a(n1688), .b(n1304), .O(n1689));
  nor2   g1374(.a(n1689), .b(n1687), .O(n1690));
  nor2   g1375(.a(G2204), .b(G18), .O(n1691));
  nor2   g1376(.a(n385), .b(n397), .O(n1692));
  nor2   g1377(.a(n1692), .b(n1691), .O(n1693));
  nor2   g1378(.a(n1693), .b(n1312), .O(n1694));
  inv1   g1379(.a(n1693), .O(n1695));
  nor2   g1380(.a(n1695), .b(n1311), .O(n1696));
  nor2   g1381(.a(n1696), .b(n1694), .O(n1697));
  inv1   g1382(.a(n1697), .O(n1698));
  nor2   g1383(.a(G114), .b(G18), .O(n1699));
  inv1   g1384(.a(G1459), .O(n1700));
  nor2   g1385(.a(n1700), .b(n397), .O(n1701));
  nor2   g1386(.a(n1701), .b(n1699), .O(n1702));
  nor2   g1387(.a(n1702), .b(n1330), .O(n1703));
  inv1   g1388(.a(n1702), .O(n1704));
  nor2   g1389(.a(n1704), .b(n1329), .O(n1705));
  nor2   g1390(.a(n1705), .b(n1703), .O(n1706));
  nor2   g1391(.a(n1706), .b(n1353), .O(n1707));
  inv1   g1392(.a(n1706), .O(n1708));
  nor2   g1393(.a(n1708), .b(n1344), .O(n1709));
  nor2   g1394(.a(n1709), .b(n1707), .O(n1710));
  inv1   g1395(.a(n1710), .O(n1711));
  nor2   g1396(.a(n1711), .b(n1698), .O(n1712));
  nor2   g1397(.a(n1710), .b(n1697), .O(n1713));
  nor2   g1398(.a(n1713), .b(n1712), .O(n1714));
  nor2   g1399(.a(n1714), .b(n1356), .O(n1715));
  inv1   g1400(.a(n1714), .O(n1716));
  nor2   g1401(.a(n1716), .b(n1349), .O(n1717));
  nor2   g1402(.a(n1717), .b(n1715), .O(n1718));
  nor2   g1403(.a(n1718), .b(n1690), .O(n1719));
  inv1   g1404(.a(n1690), .O(n1720));
  inv1   g1405(.a(n1718), .O(n1721));
  nor2   g1406(.a(n1721), .b(n1720), .O(n1722));
  nor2   g1407(.a(G3701), .b(n397), .O(n1723));
  nor2   g1408(.a(n1723), .b(n893), .O(n1724));
  inv1   g1409(.a(n1724), .O(n1725));
  nor2   g1410(.a(n888), .b(n904), .O(n1726));
  nor2   g1411(.a(n889), .b(n879), .O(n1727));
  nor2   g1412(.a(n1727), .b(n1726), .O(n1728));
  inv1   g1413(.a(n1728), .O(n1729));
  nor2   g1414(.a(n1729), .b(n1725), .O(n1730));
  nor2   g1415(.a(n1728), .b(n1724), .O(n1731));
  nor2   g1416(.a(n1731), .b(n1730), .O(n1732));
  nor2   g1417(.a(n1732), .b(n914), .O(n1733));
  inv1   g1418(.a(n1732), .O(n1734));
  nor2   g1419(.a(n1734), .b(n913), .O(n1735));
  nor2   g1420(.a(n1735), .b(n1733), .O(n1736));
  inv1   g1421(.a(n1736), .O(n1737));
  nor2   g1422(.a(n965), .b(n953), .O(n1738));
  nor2   g1423(.a(n978), .b(n945), .O(n1739));
  nor2   g1424(.a(n1739), .b(n1738), .O(n1740));
  inv1   g1425(.a(n1740), .O(n1741));
  nor2   g1426(.a(n1741), .b(n984), .O(n1742));
  nor2   g1427(.a(n1740), .b(n973), .O(n1743));
  nor2   g1428(.a(n1743), .b(n1742), .O(n1744));
  inv1   g1429(.a(n1744), .O(n1745));
  nor2   g1430(.a(G3698), .b(n397), .O(n1746));
  inv1   g1431(.a(G69), .O(n1747));
  nor2   g1432(.a(n1747), .b(G18), .O(n1748));
  nor2   g1433(.a(n1748), .b(n1746), .O(n1749));
  nor2   g1434(.a(n1749), .b(n950), .O(n1750));
  inv1   g1435(.a(n1749), .O(n1751));
  nor2   g1436(.a(n1751), .b(n937), .O(n1752));
  nor2   g1437(.a(n1752), .b(n1750), .O(n1753));
  nor2   g1438(.a(n1753), .b(n981), .O(n1754));
  inv1   g1439(.a(n1753), .O(n1755));
  nor2   g1440(.a(n1755), .b(n926), .O(n1756));
  nor2   g1441(.a(n1756), .b(n1754), .O(n1757));
  nor2   g1442(.a(n1757), .b(n1745), .O(n1758));
  inv1   g1443(.a(n1757), .O(n1759));
  nor2   g1444(.a(n1759), .b(n1744), .O(n1760));
  nor2   g1445(.a(n1760), .b(n1758), .O(n1761));
  inv1   g1446(.a(n1761), .O(n1762));
  nor2   g1447(.a(n1762), .b(n1737), .O(n1763));
  nor2   g1448(.a(n1761), .b(n1736), .O(n1764));
  nor2   g1449(.a(n1764), .b(n1763), .O(n1765));
  inv1   g1450(.a(n1765), .O(n1766));
  nor2   g1451(.a(n1766), .b(n1722), .O(n1767));
  inv1   g1452(.a(n1767), .O(n1768));
  nor2   g1453(.a(n1768), .b(n1719), .O(n1769));
  inv1   g1454(.a(n1769), .O(n1770));
  nor2   g1455(.a(n1770), .b(n1683), .O(n1771));
  inv1   g1456(.a(n1771), .O(n1772));
  nor2   g1457(.a(n1772), .b(n1680), .O(n1773));
  inv1   g1458(.a(n1773), .O(n1774));
  nor2   g1459(.a(n1774), .b(n1644), .O(n1775));
  inv1   g1460(.a(n1775), .O(G414));
  inv1   g1461(.a(n1169), .O(n1777));
  nor2   g1462(.a(n1245), .b(n1777), .O(n1778));
  inv1   g1463(.a(n1243), .O(n1779));
  nor2   g1464(.a(n1779), .b(n1171), .O(n1780));
  nor2   g1465(.a(n1780), .b(n1778), .O(n1781));
  nor2   g1466(.a(n1781), .b(n1226), .O(n1782));
  inv1   g1467(.a(n1781), .O(n1783));
  nor2   g1468(.a(n1783), .b(n1225), .O(n1784));
  nor2   g1469(.a(n1784), .b(n1782), .O(n1785));
  nor2   g1470(.a(n1785), .b(n1263), .O(n1786));
  inv1   g1471(.a(n1785), .O(n1787));
  nor2   g1472(.a(n1787), .b(n1193), .O(n1788));
  nor2   g1473(.a(n1788), .b(n1786), .O(n1789));
  inv1   g1474(.a(n1789), .O(n1790));
  inv1   g1475(.a(G181), .O(n1791));
  nor2   g1476(.a(n1791), .b(n397), .O(n1792));
  nor2   g1477(.a(n1792), .b(n1558), .O(n1793));
  inv1   g1478(.a(n1793), .O(n1794));
  inv1   g1479(.a(n1151), .O(n1795));
  nor2   g1480(.a(n1177), .b(n1795), .O(n1796));
  inv1   g1481(.a(n1159), .O(n1797));
  nor2   g1482(.a(n1797), .b(n1257), .O(n1798));
  nor2   g1483(.a(n1798), .b(n1796), .O(n1799));
  nor2   g1484(.a(n1799), .b(n1234), .O(n1800));
  inv1   g1485(.a(n1799), .O(n1801));
  nor2   g1486(.a(n1801), .b(n1211), .O(n1802));
  nor2   g1487(.a(n1802), .b(n1800), .O(n1803));
  nor2   g1488(.a(n1803), .b(n1794), .O(n1804));
  inv1   g1489(.a(n1803), .O(n1805));
  nor2   g1490(.a(n1805), .b(n1793), .O(n1806));
  nor2   g1491(.a(n1806), .b(n1804), .O(n1807));
  inv1   g1492(.a(n1807), .O(n1808));
  nor2   g1493(.a(n1808), .b(n1790), .O(n1809));
  nor2   g1494(.a(n1807), .b(n1789), .O(n1810));
  nor2   g1495(.a(n1810), .b(n1809), .O(n1811));
  nor2   g1496(.a(n1203), .b(n1185), .O(n1812));
  nor2   g1497(.a(n1266), .b(n1184), .O(n1813));
  nor2   g1498(.a(n1813), .b(n1812), .O(n1814));
  nor2   g1499(.a(n1814), .b(n1811), .O(n1815));
  inv1   g1500(.a(G197), .O(n1816));
  nor2   g1501(.a(n1816), .b(n397), .O(n1817));
  nor2   g1502(.a(n1817), .b(n1450), .O(n1818));
  nor2   g1503(.a(n1818), .b(n1064), .O(n1819));
  inv1   g1504(.a(n1818), .O(n1820));
  nor2   g1505(.a(n1820), .b(n1053), .O(n1821));
  nor2   g1506(.a(n1821), .b(n1819), .O(n1822));
  inv1   g1507(.a(n1822), .O(n1823));
  nor2   g1508(.a(n1823), .b(n1061), .O(n1824));
  nor2   g1509(.a(n1822), .b(n1032), .O(n1825));
  nor2   g1510(.a(n1825), .b(n1824), .O(n1826));
  nor2   g1511(.a(n1826), .b(n1102), .O(n1827));
  inv1   g1512(.a(n1826), .O(n1828));
  nor2   g1513(.a(n1828), .b(n1096), .O(n1829));
  nor2   g1514(.a(n1829), .b(n1827), .O(n1830));
  nor2   g1515(.a(n1112), .b(n1023), .O(n1831));
  nor2   g1516(.a(n1120), .b(n1022), .O(n1832));
  nor2   g1517(.a(n1832), .b(n1831), .O(n1833));
  nor2   g1518(.a(n1833), .b(n1087), .O(n1834));
  inv1   g1519(.a(n1833), .O(n1835));
  nor2   g1520(.a(n1835), .b(n1086), .O(n1836));
  nor2   g1521(.a(n1836), .b(n1834), .O(n1837));
  inv1   g1522(.a(n1837), .O(n1838));
  nor2   g1523(.a(n1838), .b(n1130), .O(n1839));
  nor2   g1524(.a(n1837), .b(n1129), .O(n1840));
  nor2   g1525(.a(n1840), .b(n1839), .O(n1841));
  inv1   g1526(.a(n1841), .O(n1842));
  nor2   g1527(.a(n1012), .b(n1042), .O(n1843));
  nor2   g1528(.a(n1045), .b(n1004), .O(n1844));
  nor2   g1529(.a(n1844), .b(n1843), .O(n1845));
  nor2   g1530(.a(n1845), .b(n1842), .O(n1846));
  inv1   g1531(.a(n1845), .O(n1847));
  nor2   g1532(.a(n1847), .b(n1841), .O(n1848));
  nor2   g1533(.a(n1848), .b(n1846), .O(n1849));
  nor2   g1534(.a(n1849), .b(n1830), .O(n1850));
  inv1   g1535(.a(n1811), .O(n1851));
  inv1   g1536(.a(n1814), .O(n1852));
  nor2   g1537(.a(n1852), .b(n1851), .O(n1853));
  nor2   g1538(.a(n1853), .b(n1850), .O(n1854));
  inv1   g1539(.a(n1854), .O(n1855));
  nor2   g1540(.a(n1855), .b(n1815), .O(n1856));
  inv1   g1541(.a(n1856), .O(n1857));
  nor2   g1542(.a(n980), .b(n883), .O(n1858));
  nor2   g1543(.a(n922), .b(n884), .O(n1859));
  nor2   g1544(.a(n1859), .b(n1858), .O(n1860));
  nor2   g1545(.a(n1860), .b(n977), .O(n1861));
  inv1   g1546(.a(n1860), .O(n1862));
  nor2   g1547(.a(n1862), .b(n961), .O(n1863));
  nor2   g1548(.a(n1863), .b(n1861), .O(n1864));
  inv1   g1549(.a(n1864), .O(n1865));
  inv1   g1550(.a(G208), .O(n1866));
  nor2   g1551(.a(n1866), .b(n397), .O(n1867));
  nor2   g1552(.a(n1867), .b(n1483), .O(n1868));
  inv1   g1553(.a(n1868), .O(n1869));
  inv1   g1554(.a(G198), .O(n1870));
  nor2   g1555(.a(n1870), .b(n397), .O(n1871));
  nor2   g1556(.a(n1871), .b(n373), .O(n1872));
  nor2   g1557(.a(n1872), .b(n903), .O(n1873));
  inv1   g1558(.a(n1872), .O(n1874));
  nor2   g1559(.a(n1874), .b(n875), .O(n1875));
  nor2   g1560(.a(n1875), .b(n1873), .O(n1876));
  inv1   g1561(.a(n1876), .O(n1877));
  nor2   g1562(.a(n1877), .b(n1869), .O(n1878));
  nor2   g1563(.a(n1876), .b(n1868), .O(n1879));
  nor2   g1564(.a(n1879), .b(n1878), .O(n1880));
  nor2   g1565(.a(n949), .b(n908), .O(n1881));
  nor2   g1566(.a(n933), .b(n909), .O(n1882));
  nor2   g1567(.a(n1882), .b(n1881), .O(n1883));
  inv1   g1568(.a(n1883), .O(n1884));
  nor2   g1569(.a(n1884), .b(n952), .O(n1885));
  nor2   g1570(.a(n1883), .b(n941), .O(n1886));
  nor2   g1571(.a(n1886), .b(n1885), .O(n1887));
  nor2   g1572(.a(n1887), .b(n983), .O(n1888));
  inv1   g1573(.a(n1887), .O(n1889));
  nor2   g1574(.a(n1889), .b(n969), .O(n1890));
  nor2   g1575(.a(n1890), .b(n1888), .O(n1891));
  inv1   g1576(.a(n1891), .O(n1892));
  nor2   g1577(.a(n1892), .b(n1880), .O(n1893));
  inv1   g1578(.a(n1880), .O(n1894));
  nor2   g1579(.a(n1891), .b(n1894), .O(n1895));
  nor2   g1580(.a(n1895), .b(n1893), .O(n1896));
  nor2   g1581(.a(n1896), .b(n1865), .O(n1897));
  inv1   g1582(.a(n1896), .O(n1898));
  nor2   g1583(.a(n1898), .b(n1864), .O(n1899));
  nor2   g1584(.a(n1899), .b(n1897), .O(n1900));
  inv1   g1585(.a(n1830), .O(n1901));
  inv1   g1586(.a(n1849), .O(n1902));
  nor2   g1587(.a(n1902), .b(n1901), .O(n1903));
  inv1   g1588(.a(n1306), .O(n1904));
  inv1   g1589(.a(n1338), .O(n1905));
  nor2   g1590(.a(G170), .b(n397), .O(n1906));
  nor2   g1591(.a(n1906), .b(n1298), .O(n1907));
  inv1   g1592(.a(n1298), .O(n1908));
  inv1   g1593(.a(n1906), .O(n1909));
  nor2   g1594(.a(n1909), .b(n1908), .O(n1910));
  nor2   g1595(.a(n1910), .b(n1907), .O(n1911));
  inv1   g1596(.a(n1911), .O(n1912));
  nor2   g1597(.a(n1912), .b(n1905), .O(n1913));
  nor2   g1598(.a(n1911), .b(n1338), .O(n1914));
  nor2   g1599(.a(n1914), .b(n1913), .O(n1915));
  nor2   g1600(.a(n1915), .b(n1324), .O(n1916));
  inv1   g1601(.a(n1324), .O(n1917));
  inv1   g1602(.a(n1915), .O(n1918));
  nor2   g1603(.a(n1918), .b(n1917), .O(n1919));
  nor2   g1604(.a(n1919), .b(n1916), .O(n1920));
  inv1   g1605(.a(n1920), .O(n1921));
  nor2   g1606(.a(n1921), .b(n1904), .O(n1922));
  nor2   g1607(.a(n1920), .b(n1306), .O(n1923));
  nor2   g1608(.a(n1923), .b(n1922), .O(n1924));
  inv1   g1609(.a(n1924), .O(n1925));
  inv1   g1610(.a(G164), .O(n1926));
  nor2   g1611(.a(G165), .b(n1926), .O(n1927));
  inv1   g1612(.a(G165), .O(n1928));
  nor2   g1613(.a(n1928), .b(G164), .O(n1929));
  nor2   g1614(.a(n1929), .b(n1927), .O(n1930));
  nor2   g1615(.a(n1930), .b(n1521), .O(n1931));
  nor2   g1616(.a(n1931), .b(n396), .O(n1932));
  inv1   g1617(.a(n1932), .O(n1933));
  nor2   g1618(.a(n1933), .b(n1925), .O(n1934));
  inv1   g1619(.a(n1931), .O(n1935));
  nor2   g1620(.a(n1935), .b(n1924), .O(n1936));
  nor2   g1621(.a(n1936), .b(n1934), .O(n1937));
  inv1   g1622(.a(n1937), .O(n1938));
  nor2   g1623(.a(n1938), .b(n1903), .O(n1939));
  inv1   g1624(.a(n1939), .O(n1940));
  nor2   g1625(.a(n1940), .b(n1900), .O(n1941));
  inv1   g1626(.a(n1941), .O(n1942));
  nor2   g1627(.a(n1942), .b(n1857), .O(n1943));
  inv1   g1628(.a(n1943), .O(G416));
  nor2   g1629(.a(n759), .b(n713), .O(n1945));
  inv1   g1630(.a(n713), .O(n1946));
  nor2   g1631(.a(n758), .b(n1946), .O(n1947));
  nor2   g1632(.a(n1947), .b(n1945), .O(G295));
  nor2   g1633(.a(n813), .b(n797), .O(n1949));
  inv1   g1634(.a(n797), .O(n1950));
  nor2   g1635(.a(n812), .b(n1950), .O(n1951));
  nor2   g1636(.a(n1951), .b(n1949), .O(G324));
  inv1   g1637(.a(n1150), .O(G252));
  nor2   g1638(.a(n784), .b(n762), .O(n1954));
  nor2   g1639(.a(n784), .b(n1946), .O(n1955));
  nor2   g1640(.a(n1955), .b(n1954), .O(n1956));
  nor2   g1641(.a(n1956), .b(n771), .O(n1957));
  inv1   g1642(.a(n1956), .O(n1958));
  nor2   g1643(.a(n1958), .b(n770), .O(n1959));
  nor2   g1644(.a(n1959), .b(n1957), .O(n1960));
  inv1   g1645(.a(n1960), .O(G310));
  inv1   g1646(.a(n781), .O(n1962));
  nor2   g1647(.a(n1962), .b(n1946), .O(n1963));
  inv1   g1648(.a(n779), .O(n1964));
  nor2   g1649(.a(n1964), .b(n760), .O(n1965));
  nor2   g1650(.a(n1965), .b(n733), .O(n1966));
  nor2   g1651(.a(n1966), .b(n730), .O(n1967));
  nor2   g1652(.a(n1967), .b(n1963), .O(n1968));
  inv1   g1653(.a(n1968), .O(n1969));
  nor2   g1654(.a(n1969), .b(n723), .O(n1970));
  nor2   g1655(.a(n1968), .b(n724), .O(n1971));
  nor2   g1656(.a(n1971), .b(n1970), .O(n1972));
  inv1   g1657(.a(n1972), .O(G313));
  nor2   g1658(.a(n1945), .b(n754), .O(n1974));
  nor2   g1659(.a(n1974), .b(n748), .O(n1975));
  nor2   g1660(.a(n1975), .b(n743), .O(n1976));
  inv1   g1661(.a(n1976), .O(n1977));
  nor2   g1662(.a(n1977), .b(n734), .O(n1978));
  nor2   g1663(.a(n1976), .b(n735), .O(n1979));
  nor2   g1664(.a(n1979), .b(n1978), .O(G316));
  inv1   g1665(.a(n1974), .O(n1981));
  nor2   g1666(.a(n1981), .b(n747), .O(n1982));
  nor2   g1667(.a(n1982), .b(n1975), .O(G319));
  nor2   g1668(.a(n815), .b(n797), .O(n1984));
  inv1   g1669(.a(n1984), .O(n1985));
  nor2   g1670(.a(n1985), .b(n833), .O(n1986));
  nor2   g1671(.a(n1986), .b(n854), .O(n1987));
  inv1   g1672(.a(n1987), .O(n1988));
  nor2   g1673(.a(n1988), .b(n843), .O(n1989));
  nor2   g1674(.a(n1987), .b(n842), .O(n1990));
  nor2   g1675(.a(n1990), .b(n1989), .O(n1991));
  inv1   g1676(.a(n1991), .O(G327));
  nor2   g1677(.a(n1984), .b(n850), .O(n1993));
  nor2   g1678(.a(n1993), .b(n829), .O(n1994));
  nor2   g1679(.a(n1994), .b(n827), .O(n1995));
  nor2   g1680(.a(n1995), .b(n823), .O(n1996));
  inv1   g1681(.a(n1995), .O(n1997));
  nor2   g1682(.a(n1997), .b(n822), .O(n1998));
  nor2   g1683(.a(n1998), .b(n1996), .O(G330));
  nor2   g1684(.a(n1993), .b(n831), .O(n2000));
  inv1   g1685(.a(n1993), .O(n2001));
  nor2   g1686(.a(n2001), .b(n830), .O(n2002));
  nor2   g1687(.a(n2002), .b(n2000), .O(G333));
  nor2   g1688(.a(n809), .b(n804), .O(n2004));
  nor2   g1689(.a(n2004), .b(n848), .O(n2005));
  nor2   g1690(.a(n2005), .b(n1949), .O(n2006));
  nor2   g1691(.a(n2006), .b(n1984), .O(G336));
  nor2   g1692(.a(G406), .b(G404), .O(n2008));
  inv1   g1693(.a(n2008), .O(n2009));
  nor2   g1694(.a(G410), .b(G408), .O(n2010));
  inv1   g1695(.a(n2010), .O(n2011));
  nor2   g1696(.a(n2011), .b(n2009), .O(n2012));
  inv1   g1697(.a(n2012), .O(n2013));
  nor2   g1698(.a(n2013), .b(G416), .O(n2014));
  inv1   g1699(.a(n2014), .O(n2015));
  nor2   g1700(.a(n2015), .b(G412), .O(n2016));
  inv1   g1701(.a(n2016), .O(n2017));
  nor2   g1702(.a(n2017), .b(G414), .O(n2018));
  inv1   g1703(.a(n2018), .O(G418));
  nor2   g1704(.a(n786), .b(n774), .O(n2020));
  nor2   g1705(.a(n2020), .b(n437), .O(n2021));
  nor2   g1706(.a(n2021), .b(n790), .O(n2022));
  nor2   g1707(.a(n2022), .b(n405), .O(n2023));
  inv1   g1708(.a(n2022), .O(n2024));
  nor2   g1709(.a(n2024), .b(n404), .O(n2025));
  nor2   g1710(.a(n2025), .b(n2023), .O(G298));
  nor2   g1711(.a(n429), .b(n409), .O(n2027));
  inv1   g1712(.a(n2027), .O(n2028));
  inv1   g1713(.a(n2020), .O(n2029));
  nor2   g1714(.a(n2029), .b(n425), .O(n2030));
  nor2   g1715(.a(n2030), .b(n433), .O(n2031));
  nor2   g1716(.a(n2031), .b(n2028), .O(n2032));
  inv1   g1717(.a(n2031), .O(n2033));
  nor2   g1718(.a(n2033), .b(n2027), .O(n2034));
  nor2   g1719(.a(n2034), .b(n2032), .O(n2035));
  inv1   g1720(.a(n2035), .O(G301));
  nor2   g1721(.a(n431), .b(n421), .O(n2037));
  inv1   g1722(.a(n2037), .O(n2038));
  nor2   g1723(.a(n2038), .b(n2029), .O(n2039));
  inv1   g1724(.a(n431), .O(n2040));
  nor2   g1725(.a(n2040), .b(n416), .O(n2041));
  nor2   g1726(.a(n2041), .b(n432), .O(n2042));
  inv1   g1727(.a(n2042), .O(n2043));
  nor2   g1728(.a(n2043), .b(n2039), .O(n2044));
  inv1   g1729(.a(n2039), .O(n2045));
  nor2   g1730(.a(n2045), .b(n417), .O(n2046));
  nor2   g1731(.a(n2046), .b(n2044), .O(n2047));
  inv1   g1732(.a(n2047), .O(G304));
  nor2   g1733(.a(n2037), .b(n2020), .O(n2049));
  nor2   g1734(.a(n2049), .b(n2039), .O(n2050));
  inv1   g1735(.a(n2050), .O(G307));
  nor2   g1736(.a(n1412), .b(n489), .O(n2052));
  nor2   g1737(.a(n2052), .b(n549), .O(n2053));
  nor2   g1738(.a(n2053), .b(n650), .O(n2054));
  inv1   g1739(.a(n2053), .O(n2055));
  nor2   g1740(.a(n2055), .b(n649), .O(n2056));
  nor2   g1741(.a(n2056), .b(n2054), .O(G344));
  inv1   g1742(.a(n389), .O(n2058));
  nor2   g1743(.a(n2058), .b(n868), .O(n2059));
  nor2   g1744(.a(n2059), .b(n390), .O(n2060));
  nor2   g1745(.a(n2060), .b(n862), .O(n2061));
  nor2   g1746(.a(n390), .b(n863), .O(n2062));
  nor2   g1747(.a(n2062), .b(n392), .O(n2063));
  inv1   g1748(.a(n2063), .O(n2064));
  nor2   g1749(.a(n2064), .b(n2061), .O(n2065));
  inv1   g1750(.a(n2061), .O(n2066));
  nor2   g1751(.a(n2063), .b(n2066), .O(n2067));
  nor2   g1752(.a(n2067), .b(n2065), .O(n2068));
  inv1   g1753(.a(n2068), .O(G422));
  inv1   g1754(.a(n2060), .O(n2070));
  nor2   g1755(.a(n2070), .b(n859), .O(n2071));
  nor2   g1756(.a(n2071), .b(n2061), .O(n2072));
  inv1   g1757(.a(n2072), .O(G419));
  inv1   g1758(.a(n675), .O(n2074));
  nor2   g1759(.a(n678), .b(n2074), .O(n2075));
  nor2   g1760(.a(n2075), .b(n624), .O(n2076));
  nor2   g1761(.a(n2076), .b(n621), .O(n2077));
  inv1   g1762(.a(n2077), .O(n2078));
  inv1   g1763(.a(n2075), .O(n2079));
  nor2   g1764(.a(n2053), .b(n665), .O(n2080));
  nor2   g1765(.a(n2080), .b(n2079), .O(n2081));
  nor2   g1766(.a(n2081), .b(n626), .O(n2082));
  nor2   g1767(.a(n2082), .b(n2078), .O(n2083));
  inv1   g1768(.a(n2083), .O(n2084));
  nor2   g1769(.a(n2084), .b(n614), .O(n2085));
  nor2   g1770(.a(n2083), .b(n615), .O(n2086));
  nor2   g1771(.a(n2086), .b(n2085), .O(G359));
  inv1   g1772(.a(n2081), .O(n2088));
  nor2   g1773(.a(n2088), .b(n625), .O(n2089));
  nor2   g1774(.a(n2089), .b(n2082), .O(G362));
  nor2   g1775(.a(n2053), .b(n652), .O(n2091));
  nor2   g1776(.a(n2091), .b(n672), .O(n2092));
  inv1   g1777(.a(n2092), .O(n2093));
  nor2   g1778(.a(n2093), .b(n634), .O(n2094));
  nor2   g1779(.a(n2094), .b(n663), .O(n2095));
  inv1   g1780(.a(n2094), .O(n2096));
  nor2   g1781(.a(n2096), .b(n662), .O(n2097));
  nor2   g1782(.a(n2097), .b(n2095), .O(G365));
  nor2   g1783(.a(n645), .b(n638), .O(n2099));
  inv1   g1784(.a(n2099), .O(n2100));
  nor2   g1785(.a(n2100), .b(n2054), .O(n2101));
  nor2   g1786(.a(n2101), .b(n2093), .O(G368));
  inv1   g1787(.a(n2080), .O(n2103));
  nor2   g1788(.a(n2103), .b(n628), .O(n2104));
  nor2   g1789(.a(n2104), .b(n688), .O(n2105));
  nor2   g1790(.a(n2105), .b(n602), .O(n2106));
  nor2   g1791(.a(n2106), .b(n708), .O(n2107));
  inv1   g1792(.a(n2107), .O(n2108));
  nor2   g1793(.a(n2108), .b(n560), .O(n2109));
  nor2   g1794(.a(n2107), .b(n561), .O(n2110));
  nor2   g1795(.a(n2110), .b(n2109), .O(G347));
  nor2   g1796(.a(n593), .b(n569), .O(n2112));
  inv1   g1797(.a(n2112), .O(n2113));
  inv1   g1798(.a(n2105), .O(n2114));
  nor2   g1799(.a(n2114), .b(n590), .O(n2115));
  nor2   g1800(.a(n2115), .b(n598), .O(n2116));
  nor2   g1801(.a(n2116), .b(n2113), .O(n2117));
  inv1   g1802(.a(n2116), .O(n2118));
  nor2   g1803(.a(n2118), .b(n2112), .O(n2119));
  nor2   g1804(.a(n2119), .b(n2117), .O(n2120));
  inv1   g1805(.a(n2120), .O(G350));
  nor2   g1806(.a(n596), .b(n586), .O(n2122));
  inv1   g1807(.a(n2122), .O(n2123));
  nor2   g1808(.a(n2123), .b(n2114), .O(n2124));
  inv1   g1809(.a(n596), .O(n2125));
  nor2   g1810(.a(n2125), .b(n579), .O(n2126));
  nor2   g1811(.a(n2126), .b(n597), .O(n2127));
  inv1   g1812(.a(n2127), .O(n2128));
  nor2   g1813(.a(n2128), .b(n2124), .O(n2129));
  inv1   g1814(.a(n2124), .O(n2130));
  nor2   g1815(.a(n2130), .b(n580), .O(n2131));
  nor2   g1816(.a(n2131), .b(n2129), .O(n2132));
  inv1   g1817(.a(n2132), .O(G353));
  nor2   g1818(.a(n2122), .b(n2105), .O(n2134));
  nor2   g1819(.a(n2134), .b(n2124), .O(n2135));
  inv1   g1820(.a(n2135), .O(G356));
  nor2   g1821(.a(n429), .b(n424), .O(n2137));
  nor2   g1822(.a(n2137), .b(n426), .O(n2138));
  nor2   g1823(.a(n2138), .b(n405), .O(n2139));
  inv1   g1824(.a(n2138), .O(n2140));
  nor2   g1825(.a(n2140), .b(n404), .O(n2141));
  nor2   g1826(.a(n2141), .b(n2139), .O(n2142));
  inv1   g1827(.a(n2142), .O(n2143));
  nor2   g1828(.a(n2143), .b(n2043), .O(n2144));
  nor2   g1829(.a(n2142), .b(n2042), .O(n2145));
  nor2   g1830(.a(n2145), .b(n2144), .O(n2146));
  inv1   g1831(.a(n2146), .O(n2147));
  nor2   g1832(.a(n2147), .b(n2029), .O(n2148));
  inv1   g1833(.a(n433), .O(n2149));
  nor2   g1834(.a(n2149), .b(n409), .O(n2150));
  nor2   g1835(.a(n2150), .b(n434), .O(n2151));
  inv1   g1836(.a(n2151), .O(n2152));
  nor2   g1837(.a(n421), .b(n416), .O(n2153));
  nor2   g1838(.a(n2153), .b(n423), .O(n2154));
  nor2   g1839(.a(n2154), .b(n405), .O(n2155));
  inv1   g1840(.a(n2154), .O(n2156));
  nor2   g1841(.a(n2156), .b(n404), .O(n2157));
  nor2   g1842(.a(n2157), .b(n2155), .O(n2158));
  nor2   g1843(.a(n2158), .b(n2152), .O(n2159));
  inv1   g1844(.a(n2158), .O(n2160));
  nor2   g1845(.a(n2160), .b(n2151), .O(n2161));
  nor2   g1846(.a(n2161), .b(n2159), .O(n2162));
  inv1   g1847(.a(n2162), .O(n2163));
  nor2   g1848(.a(n2163), .b(n2020), .O(n2164));
  nor2   g1849(.a(n2164), .b(n2148), .O(n2165));
  inv1   g1850(.a(n2165), .O(n2166));
  nor2   g1851(.a(n1964), .b(n730), .O(n2167));
  nor2   g1852(.a(n2167), .b(n780), .O(n2168));
  inv1   g1853(.a(n2168), .O(n2169));
  nor2   g1854(.a(n2169), .b(n723), .O(n2170));
  nor2   g1855(.a(n734), .b(n723), .O(n2171));
  nor2   g1856(.a(n2171), .b(n736), .O(n2172));
  inv1   g1857(.a(n2172), .O(n2173));
  nor2   g1858(.a(n2173), .b(n2168), .O(n2174));
  nor2   g1859(.a(n2174), .b(n2170), .O(n2175));
  inv1   g1860(.a(n2175), .O(n2176));
  inv1   g1861(.a(n757), .O(n2177));
  nor2   g1862(.a(n770), .b(n748), .O(n2178));
  nor2   g1863(.a(n771), .b(n747), .O(n2179));
  nor2   g1864(.a(n2179), .b(n2178), .O(n2180));
  inv1   g1865(.a(n2180), .O(n2181));
  nor2   g1866(.a(n2181), .b(n2177), .O(n2182));
  nor2   g1867(.a(n2180), .b(n757), .O(n2183));
  nor2   g1868(.a(n2183), .b(n2182), .O(n2184));
  nor2   g1869(.a(n2184), .b(n784), .O(n2185));
  inv1   g1870(.a(n2184), .O(n2186));
  nor2   g1871(.a(n2186), .b(n783), .O(n2187));
  nor2   g1872(.a(n2187), .b(n2185), .O(n2188));
  nor2   g1873(.a(n2188), .b(n2176), .O(n2189));
  inv1   g1874(.a(n2188), .O(n2190));
  nor2   g1875(.a(n2190), .b(n2175), .O(n2191));
  nor2   g1876(.a(n2191), .b(n2189), .O(n2192));
  nor2   g1877(.a(n2192), .b(n1946), .O(n2193));
  inv1   g1878(.a(n1967), .O(n2194));
  nor2   g1879(.a(n2180), .b(n2194), .O(n2195));
  nor2   g1880(.a(n2181), .b(n1967), .O(n2196));
  nor2   g1881(.a(n2196), .b(n2195), .O(n2197));
  inv1   g1882(.a(n2197), .O(n2198));
  inv1   g1883(.a(n1965), .O(n2199));
  nor2   g1884(.a(n2199), .b(n783), .O(n2200));
  inv1   g1885(.a(n1954), .O(n2201));
  nor2   g1886(.a(n1965), .b(n2201), .O(n2202));
  nor2   g1887(.a(n2202), .b(n2200), .O(n2203));
  inv1   g1888(.a(n2203), .O(n2204));
  nor2   g1889(.a(n2172), .b(n777), .O(n2205));
  nor2   g1890(.a(n2173), .b(n754), .O(n2206));
  nor2   g1891(.a(n2206), .b(n2205), .O(n2207));
  nor2   g1892(.a(n2207), .b(n2204), .O(n2208));
  inv1   g1893(.a(n2207), .O(n2209));
  nor2   g1894(.a(n2209), .b(n2203), .O(n2210));
  nor2   g1895(.a(n2210), .b(n2208), .O(n2211));
  nor2   g1896(.a(n2211), .b(n2198), .O(n2212));
  inv1   g1897(.a(n2211), .O(n2213));
  nor2   g1898(.a(n2213), .b(n2197), .O(n2214));
  nor2   g1899(.a(n2214), .b(n2212), .O(n2215));
  nor2   g1900(.a(n2215), .b(n713), .O(n2216));
  nor2   g1901(.a(n2216), .b(n2193), .O(n2217));
  nor2   g1902(.a(n2217), .b(n2166), .O(n2218));
  inv1   g1903(.a(n2217), .O(n2219));
  nor2   g1904(.a(n2219), .b(n2165), .O(n2220));
  nor2   g1905(.a(n2220), .b(n2218), .O(n2221));
  inv1   g1906(.a(n2221), .O(G321));
  nor2   g1907(.a(n2063), .b(n862), .O(n2223));
  inv1   g1908(.a(n2059), .O(n2224));
  nor2   g1909(.a(n2224), .b(G1496), .O(n2225));
  nor2   g1910(.a(n2059), .b(n863), .O(n2226));
  nor2   g1911(.a(n2226), .b(n2225), .O(n2227));
  inv1   g1912(.a(n2227), .O(n2228));
  nor2   g1913(.a(n2228), .b(n859), .O(n2229));
  nor2   g1914(.a(n2229), .b(n2223), .O(n2230));
  inv1   g1915(.a(n2230), .O(n2231));
  nor2   g1916(.a(n848), .b(n803), .O(n2232));
  inv1   g1917(.a(n2232), .O(n2233));
  nor2   g1918(.a(n852), .b(n847), .O(n2234));
  nor2   g1919(.a(n827), .b(n801), .O(n2235));
  nor2   g1920(.a(n2235), .b(n829), .O(n2236));
  inv1   g1921(.a(n2236), .O(n2237));
  nor2   g1922(.a(n2237), .b(n809), .O(n2238));
  nor2   g1923(.a(n2238), .b(n812), .O(n2239));
  inv1   g1924(.a(n2239), .O(n2240));
  nor2   g1925(.a(n2240), .b(n2234), .O(n2241));
  nor2   g1926(.a(n2237), .b(n813), .O(n2242));
  nor2   g1927(.a(n2242), .b(n2241), .O(n2243));
  nor2   g1928(.a(n2243), .b(n855), .O(n2244));
  inv1   g1929(.a(n2243), .O(n2245));
  nor2   g1930(.a(n2245), .b(n854), .O(n2246));
  nor2   g1931(.a(n2246), .b(n2244), .O(n2247));
  nor2   g1932(.a(n830), .b(n822), .O(n2248));
  nor2   g1933(.a(n2248), .b(n832), .O(n2249));
  inv1   g1934(.a(n2249), .O(n2250));
  nor2   g1935(.a(n2250), .b(n843), .O(n2251));
  nor2   g1936(.a(n2249), .b(n842), .O(n2252));
  nor2   g1937(.a(n2252), .b(n2251), .O(n2253));
  inv1   g1938(.a(n2253), .O(n2254));
  nor2   g1939(.a(n2254), .b(n2247), .O(n2255));
  inv1   g1940(.a(n2247), .O(n2256));
  nor2   g1941(.a(n2253), .b(n2256), .O(n2257));
  nor2   g1942(.a(n2257), .b(n2255), .O(n2258));
  inv1   g1943(.a(n2258), .O(n2259));
  nor2   g1944(.a(n2259), .b(n2233), .O(n2260));
  nor2   g1945(.a(n2258), .b(n2232), .O(n2261));
  nor2   g1946(.a(n2261), .b(n2260), .O(n2262));
  nor2   g1947(.a(n2262), .b(n1950), .O(n2263));
  nor2   g1948(.a(n854), .b(n834), .O(n2264));
  inv1   g1949(.a(n2264), .O(n2265));
  inv1   g1950(.a(n2005), .O(n2266));
  nor2   g1951(.a(n2253), .b(n2266), .O(n2267));
  nor2   g1952(.a(n2254), .b(n2005), .O(n2268));
  nor2   g1953(.a(n2268), .b(n2267), .O(n2269));
  inv1   g1954(.a(n2269), .O(n2270));
  nor2   g1955(.a(n2270), .b(n2265), .O(n2271));
  nor2   g1956(.a(n2269), .b(n2264), .O(n2272));
  nor2   g1957(.a(n2272), .b(n2271), .O(n2273));
  inv1   g1958(.a(n2273), .O(n2274));
  nor2   g1959(.a(n850), .b(n814), .O(n2275));
  nor2   g1960(.a(n2275), .b(n829), .O(n2276));
  inv1   g1961(.a(n2275), .O(n2277));
  nor2   g1962(.a(n2277), .b(n827), .O(n2278));
  nor2   g1963(.a(n2278), .b(n2276), .O(n2279));
  nor2   g1964(.a(n2279), .b(n2274), .O(n2280));
  inv1   g1965(.a(n2279), .O(n2281));
  nor2   g1966(.a(n2281), .b(n2273), .O(n2282));
  nor2   g1967(.a(n2282), .b(n2280), .O(n2283));
  nor2   g1968(.a(n2283), .b(n797), .O(n2284));
  nor2   g1969(.a(n2284), .b(n2263), .O(n2285));
  nor2   g1970(.a(n2285), .b(n2231), .O(n2286));
  inv1   g1971(.a(n2285), .O(n2287));
  nor2   g1972(.a(n2287), .b(n2230), .O(n2288));
  nor2   g1973(.a(n2288), .b(n2286), .O(G338));
  nor2   g1974(.a(n593), .b(n589), .O(n2290));
  nor2   g1975(.a(n2290), .b(n591), .O(n2291));
  nor2   g1976(.a(n2291), .b(n561), .O(n2292));
  inv1   g1977(.a(n2291), .O(n2293));
  nor2   g1978(.a(n2293), .b(n560), .O(n2294));
  nor2   g1979(.a(n2294), .b(n2292), .O(n2295));
  inv1   g1980(.a(n2295), .O(n2296));
  nor2   g1981(.a(n2296), .b(n2128), .O(n2297));
  nor2   g1982(.a(n2295), .b(n2127), .O(n2298));
  nor2   g1983(.a(n2298), .b(n2297), .O(n2299));
  inv1   g1984(.a(n2299), .O(n2300));
  nor2   g1985(.a(n2300), .b(n2114), .O(n2301));
  nor2   g1986(.a(n586), .b(n579), .O(n2302));
  nor2   g1987(.a(n2302), .b(n588), .O(n2303));
  nor2   g1988(.a(n2303), .b(n561), .O(n2304));
  inv1   g1989(.a(n2303), .O(n2305));
  nor2   g1990(.a(n2305), .b(n560), .O(n2306));
  nor2   g1991(.a(n2306), .b(n2304), .O(n2307));
  inv1   g1992(.a(n2307), .O(n2308));
  inv1   g1993(.a(n598), .O(n2309));
  nor2   g1994(.a(n2309), .b(n569), .O(n2310));
  nor2   g1995(.a(n2310), .b(n599), .O(n2311));
  nor2   g1996(.a(n2311), .b(n2308), .O(n2312));
  inv1   g1997(.a(n2311), .O(n2313));
  nor2   g1998(.a(n2313), .b(n2307), .O(n2314));
  nor2   g1999(.a(n2314), .b(n2312), .O(n2315));
  inv1   g2000(.a(n2315), .O(n2316));
  nor2   g2001(.a(n2316), .b(n2105), .O(n2317));
  nor2   g2002(.a(n2317), .b(n2301), .O(n2318));
  inv1   g2003(.a(n2318), .O(n2319));
  inv1   g2004(.a(n648), .O(n2320));
  nor2   g2005(.a(n2079), .b(n621), .O(n2321));
  nor2   g2006(.a(n2321), .b(n2076), .O(n2322));
  nor2   g2007(.a(n2322), .b(n2320), .O(n2323));
  inv1   g2008(.a(n2322), .O(n2324));
  nor2   g2009(.a(n2324), .b(n648), .O(n2325));
  nor2   g2010(.a(n2325), .b(n2323), .O(n2326));
  inv1   g2011(.a(n2326), .O(n2327));
  nor2   g2012(.a(n625), .b(n614), .O(n2328));
  nor2   g2013(.a(n2328), .b(n627), .O(n2329));
  nor2   g2014(.a(n2329), .b(n663), .O(n2330));
  inv1   g2015(.a(n2329), .O(n2331));
  nor2   g2016(.a(n2331), .b(n662), .O(n2332));
  nor2   g2017(.a(n2332), .b(n2330), .O(n2333));
  inv1   g2018(.a(n2333), .O(n2334));
  nor2   g2019(.a(n672), .b(n637), .O(n2335));
  nor2   g2020(.a(n2335), .b(n2334), .O(n2336));
  inv1   g2021(.a(n2335), .O(n2337));
  nor2   g2022(.a(n2337), .b(n2333), .O(n2338));
  nor2   g2023(.a(n2338), .b(n2336), .O(n2339));
  nor2   g2024(.a(n2339), .b(n2327), .O(n2340));
  inv1   g2025(.a(n2339), .O(n2341));
  nor2   g2026(.a(n2341), .b(n2326), .O(n2342));
  nor2   g2027(.a(n2342), .b(n2340), .O(n2343));
  nor2   g2028(.a(n2343), .b(n2055), .O(n2344));
  nor2   g2029(.a(n2099), .b(n672), .O(n2345));
  nor2   g2030(.a(n2345), .b(n2334), .O(n2346));
  inv1   g2031(.a(n2345), .O(n2347));
  nor2   g2032(.a(n2347), .b(n2333), .O(n2348));
  nor2   g2033(.a(n2348), .b(n2346), .O(n2349));
  inv1   g2034(.a(n2349), .O(n2350));
  nor2   g2035(.a(n665), .b(n624), .O(n2351));
  nor2   g2036(.a(n2351), .b(n2078), .O(n2352));
  inv1   g2037(.a(n2352), .O(n2353));
  nor2   g2038(.a(n651), .b(n634), .O(n2354));
  inv1   g2039(.a(n2354), .O(n2355));
  nor2   g2040(.a(n2355), .b(n672), .O(n2356));
  inv1   g2041(.a(n2356), .O(n2357));
  nor2   g2042(.a(n2357), .b(n2075), .O(n2358));
  nor2   g2043(.a(n2356), .b(n664), .O(n2359));
  inv1   g2044(.a(n2359), .O(n2360));
  nor2   g2045(.a(n2360), .b(n2079), .O(n2361));
  nor2   g2046(.a(n2361), .b(n2358), .O(n2362));
  nor2   g2047(.a(n2362), .b(n2353), .O(n2363));
  inv1   g2048(.a(n2362), .O(n2364));
  nor2   g2049(.a(n2364), .b(n2352), .O(n2365));
  nor2   g2050(.a(n2365), .b(n2363), .O(n2366));
  nor2   g2051(.a(n2366), .b(n2350), .O(n2367));
  inv1   g2052(.a(n2366), .O(n2368));
  nor2   g2053(.a(n2368), .b(n2349), .O(n2369));
  nor2   g2054(.a(n2369), .b(n2367), .O(n2370));
  nor2   g2055(.a(n2370), .b(n2053), .O(n2371));
  nor2   g2056(.a(n2371), .b(n2344), .O(n2372));
  nor2   g2057(.a(n2372), .b(n2319), .O(n2373));
  inv1   g2058(.a(n2372), .O(n2374));
  nor2   g2059(.a(n2374), .b(n2318), .O(n2375));
  nor2   g2060(.a(n2375), .b(n2373), .O(G370));
  nor2   g2061(.a(n1410), .b(n483), .O(n2377));
  nor2   g2062(.a(n2377), .b(n480), .O(n2378));
  inv1   g2063(.a(n2378), .O(n2379));
  inv1   g2064(.a(n448), .O(n2380));
  nor2   g2065(.a(n456), .b(n2380), .O(n2381));
  nor2   g2066(.a(n544), .b(n448), .O(n2382));
  nor2   g2067(.a(n2382), .b(n2381), .O(n2383));
  inv1   g2068(.a(n2383), .O(n2384));
  nor2   g2069(.a(n474), .b(n460), .O(n2385));
  nor2   g2070(.a(n473), .b(n461), .O(n2386));
  nor2   g2071(.a(n2386), .b(n2385), .O(n2387));
  inv1   g2072(.a(n2387), .O(n2388));
  nor2   g2073(.a(n2388), .b(n2384), .O(n2389));
  nor2   g2074(.a(n2387), .b(n2383), .O(n2390));
  nor2   g2075(.a(n2390), .b(n2389), .O(n2391));
  nor2   g2076(.a(n2391), .b(n2379), .O(n2392));
  inv1   g2077(.a(n2391), .O(n2393));
  nor2   g2078(.a(n2393), .b(n2378), .O(n2394));
  nor2   g2079(.a(n2394), .b(n2392), .O(n2395));
  nor2   g2080(.a(n2395), .b(n1429), .O(n2396));
  nor2   g2081(.a(n1426), .b(n544), .O(n2397));
  nor2   g2082(.a(n1410), .b(n462), .O(n2398));
  inv1   g2083(.a(n2398), .O(n2399));
  nor2   g2084(.a(n2399), .b(n1425), .O(n2400));
  nor2   g2085(.a(n2400), .b(n2397), .O(n2401));
  nor2   g2086(.a(n2398), .b(n480), .O(n2402));
  nor2   g2087(.a(n482), .b(n481), .O(n2403));
  nor2   g2088(.a(n2403), .b(n2402), .O(n2404));
  nor2   g2089(.a(n2404), .b(n474), .O(n2405));
  inv1   g2090(.a(n2404), .O(n2406));
  nor2   g2091(.a(n2406), .b(n473), .O(n2407));
  nor2   g2092(.a(n2407), .b(n2405), .O(n2408));
  nor2   g2093(.a(n2408), .b(n2401), .O(n2409));
  inv1   g2094(.a(n2401), .O(n2410));
  inv1   g2095(.a(n2408), .O(n2411));
  nor2   g2096(.a(n2411), .b(n2410), .O(n2412));
  nor2   g2097(.a(n2412), .b(n2409), .O(n2413));
  nor2   g2098(.a(n2413), .b(n1412), .O(n2414));
  nor2   g2099(.a(n2414), .b(n2396), .O(n2415));
  inv1   g2100(.a(n2415), .O(n2416));
  nor2   g2101(.a(n691), .b(n533), .O(n2417));
  nor2   g2102(.a(n2417), .b(n521), .O(n2418));
  nor2   g2103(.a(n535), .b(n506), .O(n2419));
  inv1   g2104(.a(n2419), .O(n2420));
  nor2   g2105(.a(n2420), .b(n2418), .O(n2421));
  nor2   g2106(.a(n2421), .b(n509), .O(n2422));
  inv1   g2107(.a(n2422), .O(n2423));
  inv1   g2108(.a(n2417), .O(n2424));
  nor2   g2109(.a(n2424), .b(n522), .O(n2425));
  nor2   g2110(.a(n2425), .b(n2418), .O(n2426));
  nor2   g2111(.a(n2426), .b(n2423), .O(n2427));
  inv1   g2112(.a(n2426), .O(n2428));
  nor2   g2113(.a(n2428), .b(n2422), .O(n2429));
  nor2   g2114(.a(n2429), .b(n2427), .O(n2430));
  nor2   g2115(.a(n499), .b(n381), .O(n2431));
  nor2   g2116(.a(n500), .b(n380), .O(n2432));
  nor2   g2117(.a(n2432), .b(n2431), .O(n2433));
  inv1   g2118(.a(n2433), .O(n2434));
  nor2   g2119(.a(n2434), .b(n694), .O(n2435));
  nor2   g2120(.a(n2433), .b(n693), .O(n2436));
  nor2   g2121(.a(n2436), .b(n2435), .O(n2437));
  inv1   g2122(.a(n2437), .O(n2438));
  inv1   g2123(.a(n379), .O(n2439));
  nor2   g2124(.a(n689), .b(n2439), .O(n2440));
  nor2   g2125(.a(n690), .b(n379), .O(n2441));
  nor2   g2126(.a(n2441), .b(n2440), .O(n2442));
  nor2   g2127(.a(n2442), .b(n2438), .O(n2443));
  inv1   g2128(.a(n2442), .O(n2444));
  nor2   g2129(.a(n2444), .b(n2437), .O(n2445));
  nor2   g2130(.a(n2445), .b(n2443), .O(n2446));
  inv1   g2131(.a(n2446), .O(n2447));
  nor2   g2132(.a(n2447), .b(n2430), .O(n2448));
  inv1   g2133(.a(n2430), .O(n2449));
  nor2   g2134(.a(n2446), .b(n2449), .O(n2450));
  nor2   g2135(.a(n2450), .b(n371), .O(n2451));
  inv1   g2136(.a(n2451), .O(n2452));
  nor2   g2137(.a(n2452), .b(n2448), .O(n2453));
  inv1   g2138(.a(n375), .O(n2454));
  inv1   g2139(.a(n531), .O(n2455));
  nor2   g2140(.a(n2455), .b(n2454), .O(n2456));
  inv1   g2141(.a(n530), .O(n2457));
  nor2   g2142(.a(n2457), .b(n375), .O(n2458));
  nor2   g2143(.a(n2458), .b(n2456), .O(n2459));
  nor2   g2144(.a(n536), .b(n509), .O(n2460));
  nor2   g2145(.a(n2460), .b(n2419), .O(n2461));
  inv1   g2146(.a(n2461), .O(n2462));
  nor2   g2147(.a(n2462), .b(n2437), .O(n2463));
  nor2   g2148(.a(n2461), .b(n2438), .O(n2464));
  nor2   g2149(.a(n2464), .b(n2463), .O(n2465));
  inv1   g2150(.a(n2465), .O(n2466));
  nor2   g2151(.a(n2466), .b(n2459), .O(n2467));
  inv1   g2152(.a(n2459), .O(n2468));
  nor2   g2153(.a(n2465), .b(n2468), .O(n2469));
  nor2   g2154(.a(n2469), .b(G4526), .O(n2470));
  inv1   g2155(.a(n2470), .O(n2471));
  nor2   g2156(.a(n2471), .b(n2467), .O(n2472));
  nor2   g2157(.a(n2472), .b(n2453), .O(n2473));
  nor2   g2158(.a(n2473), .b(n511), .O(n2474));
  inv1   g2159(.a(n2473), .O(n2475));
  nor2   g2160(.a(n2475), .b(n510), .O(n2476));
  nor2   g2161(.a(n2476), .b(n2474), .O(n2477));
  inv1   g2162(.a(n2477), .O(n2478));
  nor2   g2163(.a(n2478), .b(n2416), .O(n2479));
  nor2   g2164(.a(n2477), .b(n2415), .O(n2480));
  nor2   g2165(.a(n2480), .b(n2479), .O(n2481));
  inv1   g2166(.a(n2481), .O(G399));
  buffer g2167(.a(ING339 ), .O(G339));
  buffer g2168(.a(G1), .O(G2));
  buffer g2169(.a(G1), .O(G3));
  buffer g2170(.a(G1459), .O(G450));
  buffer g2171(.a(G1469), .O(G448));
  buffer g2172(.a(G1480), .O(G444));
  buffer g2173(.a(G1486), .O(G442));
  buffer g2174(.a(G1492), .O(G440));
  buffer g2175(.a(G1496), .O(G438));
  buffer g2176(.a(G2208), .O(G496));
  buffer g2177(.a(G2218), .O(G494));
  buffer g2178(.a(G2224), .O(G492));
  buffer g2179(.a(G2230), .O(G490));
  buffer g2180(.a(G2236), .O(G488));
  buffer g2181(.a(G2239), .O(G486));
  buffer g2182(.a(G2247), .O(G484));
  buffer g2183(.a(G2253), .O(G482));
  buffer g2184(.a(G2256), .O(G480));
  buffer g2185(.a(G3698), .O(G560));
  buffer g2186(.a(G3701), .O(G542));
  buffer g2187(.a(G3705), .O(G558));
  buffer g2188(.a(G3711), .O(G556));
  buffer g2189(.a(G3717), .O(G554));
  buffer g2190(.a(G3723), .O(G552));
  buffer g2191(.a(G3729), .O(G550));
  buffer g2192(.a(G3737), .O(G548));
  buffer g2193(.a(G3743), .O(G546));
  buffer g2194(.a(G3749), .O(G544));
  buffer g2195(.a(G4393), .O(G540));
  buffer g2196(.a(G4400), .O(G538));
  buffer g2197(.a(G4405), .O(G536));
  buffer g2198(.a(G4410), .O(G534));
  buffer g2199(.a(G4415), .O(G532));
  buffer g2200(.a(G4420), .O(G530));
  buffer g2201(.a(G4427), .O(G528));
  buffer g2202(.a(G4432), .O(G526));
  buffer g2203(.a(G4437), .O(G524));
  buffer g2204(.a(G1462), .O(G436));
  buffer g2205(.a(G2211), .O(G478));
  buffer g2206(.a(G4394), .O(G522));
  buffer g2207(.a(G1), .O(G432));
  buffer g2208(.a(G106), .O(G446));
  inv1   g2209(.a(G15), .O(G286));
  inv1   g2210(.a(n360), .O(G289));
  inv1   g2211(.a(G15), .O(G341));
  inv1   g2212(.a(n366), .O(G281));
  buffer g2213(.a(G1), .O(G453));
  inv1   g2214(.a(n1387), .O(G264));
  nor2   g2215(.a(n866), .b(n861), .O(G270));
  inv1   g2216(.a(n1387), .O(G249));
  nor2   g2217(.a(n866), .b(n861), .O(G276));
  nor2   g2218(.a(n866), .b(n861), .O(G273));
  inv1   g2219(.a(n2068), .O(G469));
  inv1   g2220(.a(n2072), .O(G471));
endmodule


