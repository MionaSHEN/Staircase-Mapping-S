// Benchmark "c880_blif" written by ABC on Sun Apr 14 20:04:57 2019

module c880_blif  ( 
    G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat, G51gat,
    G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat, G85gat,
    G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat, G101gat,
    G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat, G138gat,
    G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat, G165gat,
    G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat, G210gat,
    G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat, G261gat,
    G267gat, G268gat,
    G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat, G421gat,
    G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat, G767gat,
    G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat, G878gat,
    G879gat, G880gat  );
  input  G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat,
    G51gat, G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat,
    G85gat, G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat,
    G101gat, G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat,
    G138gat, G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat,
    G165gat, G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat,
    G210gat, G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat,
    G261gat, G267gat, G268gat;
  output G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat,
    G421gat, G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat,
    G767gat, G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat,
    G878gat, G879gat, G880gat;
  wire n87, n88, n89, n90, n91, n93, n94, n95, n96, n99, n100, n102, n103,
    n104, n105, n106, n107, n108, n109, n111, n112, n113, n114, n115, n116,
    n118, n119, n120, n121, n123, n124, n125, n127, n129, n130, n132, n133,
    n135, n137, n138, n139, n140, n141, n142, n143, n144, n146, n147, n148,
    n149, n150, n152, n154, n155, n156, n157, n158, n159, n160, n161, n162,
    n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
    n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
    n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n199,
    n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
    n382, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
    n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n409, n410, n411, n412, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n509, n510, n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n584, n585, n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607;
  inv1   g000(.a(G42gat), .O(n87));
  inv1   g001(.a(G29gat), .O(n88));
  inv1   g002(.a(G75gat), .O(n89));
  nor2   g003(.a(n89), .b(n88), .O(n90));
  inv1   g004(.a(n90), .O(n91));
  nor2   g005(.a(n91), .b(n87), .O(G388gat));
  inv1   g006(.a(G80gat), .O(n93));
  inv1   g007(.a(G36gat), .O(n94));
  nor2   g008(.a(n94), .b(n88), .O(n95));
  inv1   g009(.a(n95), .O(n96));
  nor2   g010(.a(n96), .b(n93), .O(G389gat));
  nor2   g011(.a(n96), .b(n87), .O(G390gat));
  inv1   g012(.a(G85gat), .O(n99));
  inv1   g013(.a(G86gat), .O(n100));
  nor2   g014(.a(n100), .b(n99), .O(G391gat));
  inv1   g015(.a(G13gat), .O(n102));
  inv1   g016(.a(G17gat), .O(n103));
  nor2   g017(.a(n103), .b(n102), .O(n104));
  inv1   g018(.a(n104), .O(n105));
  inv1   g019(.a(G1gat), .O(n106));
  inv1   g020(.a(G8gat), .O(n107));
  nor2   g021(.a(n107), .b(n106), .O(n108));
  inv1   g022(.a(n108), .O(n109));
  nor2   g023(.a(n109), .b(n105), .O(G418gat));
  inv1   g024(.a(G26gat), .O(n111));
  nor2   g025(.a(n111), .b(n106), .O(n112));
  inv1   g026(.a(n112), .O(n113));
  nor2   g027(.a(n113), .b(n105), .O(n114));
  inv1   g028(.a(n114), .O(n115));
  nor2   g029(.a(n115), .b(G390gat), .O(n116));
  inv1   g030(.a(n116), .O(G419gat));
  inv1   g031(.a(G59gat), .O(n118));
  nor2   g032(.a(n89), .b(n118), .O(n119));
  inv1   g033(.a(n119), .O(n120));
  nor2   g034(.a(n120), .b(n93), .O(n121));
  inv1   g035(.a(n121), .O(G420gat));
  nor2   g036(.a(n118), .b(n94), .O(n123));
  inv1   g037(.a(n123), .O(n124));
  nor2   g038(.a(n124), .b(n93), .O(n125));
  inv1   g039(.a(n125), .O(G421gat));
  nor2   g040(.a(n124), .b(n87), .O(n127));
  inv1   g041(.a(n127), .O(G422gat));
  inv1   g042(.a(G90gat), .O(n129));
  nor2   g043(.a(G88gat), .b(G87gat), .O(n130));
  nor2   g044(.a(n130), .b(n129), .O(G423gat));
  inv1   g045(.a(G390gat), .O(n132));
  nor2   g046(.a(n115), .b(n132), .O(n133));
  inv1   g047(.a(n133), .O(G446gat));
  inv1   g048(.a(G51gat), .O(n135));
  nor2   g049(.a(n113), .b(n135), .O(G447gat));
  inv1   g050(.a(G55gat), .O(n137));
  nor2   g051(.a(n137), .b(n102), .O(n138));
  inv1   g052(.a(n138), .O(n139));
  nor2   g053(.a(n139), .b(n109), .O(n140));
  inv1   g054(.a(n140), .O(n141));
  inv1   g055(.a(G68gat), .O(n142));
  nor2   g056(.a(n142), .b(n88), .O(n143));
  inv1   g057(.a(n143), .O(n144));
  nor2   g058(.a(n144), .b(n141), .O(G448gat));
  inv1   g059(.a(G74gat), .O(n146));
  nor2   g060(.a(n142), .b(n118), .O(n147));
  inv1   g061(.a(n147), .O(n148));
  nor2   g062(.a(n148), .b(n141), .O(n149));
  inv1   g063(.a(n149), .O(n150));
  nor2   g064(.a(n150), .b(n146), .O(G449gat));
  inv1   g065(.a(G89gat), .O(n152));
  nor2   g066(.a(n130), .b(n152), .O(G450gat));
  inv1   g067(.a(G91gat), .O(n154));
  inv1   g068(.a(G96gat), .O(n155));
  nor2   g069(.a(n155), .b(n154), .O(n156));
  nor2   g070(.a(G96gat), .b(G91gat), .O(n157));
  nor2   g071(.a(n157), .b(n156), .O(n158));
  inv1   g072(.a(n158), .O(n159));
  inv1   g073(.a(G121gat), .O(n160));
  nor2   g074(.a(G126gat), .b(n160), .O(n161));
  inv1   g075(.a(G126gat), .O(n162));
  nor2   g076(.a(n162), .b(G121gat), .O(n163));
  nor2   g077(.a(n163), .b(n161), .O(n164));
  nor2   g078(.a(n164), .b(n159), .O(n165));
  inv1   g079(.a(n164), .O(n166));
  nor2   g080(.a(n166), .b(n158), .O(n167));
  nor2   g081(.a(n167), .b(n165), .O(n168));
  inv1   g082(.a(n168), .O(n169));
  inv1   g083(.a(G135gat), .O(n170));
  inv1   g084(.a(G111gat), .O(n171));
  inv1   g085(.a(G116gat), .O(n172));
  nor2   g086(.a(n172), .b(n171), .O(n173));
  nor2   g087(.a(G116gat), .b(G111gat), .O(n174));
  nor2   g088(.a(n174), .b(n173), .O(n175));
  nor2   g089(.a(n175), .b(n170), .O(n176));
  inv1   g090(.a(n175), .O(n177));
  nor2   g091(.a(n177), .b(G135gat), .O(n178));
  nor2   g092(.a(n178), .b(n176), .O(n179));
  inv1   g093(.a(n179), .O(n180));
  inv1   g094(.a(G130gat), .O(n181));
  inv1   g095(.a(G101gat), .O(n182));
  nor2   g096(.a(G106gat), .b(n182), .O(n183));
  inv1   g097(.a(G106gat), .O(n184));
  nor2   g098(.a(n184), .b(G101gat), .O(n185));
  nor2   g099(.a(n185), .b(n183), .O(n186));
  nor2   g100(.a(n186), .b(n181), .O(n187));
  inv1   g101(.a(n186), .O(n188));
  nor2   g102(.a(n188), .b(G130gat), .O(n189));
  nor2   g103(.a(n189), .b(n187), .O(n190));
  nor2   g104(.a(n190), .b(n180), .O(n191));
  inv1   g105(.a(n190), .O(n192));
  nor2   g106(.a(n192), .b(n179), .O(n193));
  nor2   g107(.a(n193), .b(n191), .O(n194));
  inv1   g108(.a(n194), .O(n195));
  nor2   g109(.a(n195), .b(n169), .O(n196));
  nor2   g110(.a(n194), .b(n168), .O(n197));
  nor2   g111(.a(n197), .b(n196), .O(G767gat));
  inv1   g112(.a(G159gat), .O(n199));
  inv1   g113(.a(G165gat), .O(n200));
  nor2   g114(.a(n200), .b(n199), .O(n201));
  nor2   g115(.a(G165gat), .b(G159gat), .O(n202));
  nor2   g116(.a(n202), .b(n201), .O(n203));
  inv1   g117(.a(n203), .O(n204));
  inv1   g118(.a(G195gat), .O(n205));
  nor2   g119(.a(G201gat), .b(n205), .O(n206));
  inv1   g120(.a(G201gat), .O(n207));
  nor2   g121(.a(n207), .b(G195gat), .O(n208));
  nor2   g122(.a(n208), .b(n206), .O(n209));
  nor2   g123(.a(n209), .b(n204), .O(n210));
  inv1   g124(.a(n209), .O(n211));
  nor2   g125(.a(n211), .b(n203), .O(n212));
  nor2   g126(.a(n212), .b(n210), .O(n213));
  inv1   g127(.a(n213), .O(n214));
  inv1   g128(.a(G207gat), .O(n215));
  inv1   g129(.a(G183gat), .O(n216));
  inv1   g130(.a(G189gat), .O(n217));
  nor2   g131(.a(n217), .b(n216), .O(n218));
  nor2   g132(.a(G189gat), .b(G183gat), .O(n219));
  nor2   g133(.a(n219), .b(n218), .O(n220));
  nor2   g134(.a(n220), .b(n215), .O(n221));
  inv1   g135(.a(n220), .O(n222));
  nor2   g136(.a(n222), .b(G207gat), .O(n223));
  nor2   g137(.a(n223), .b(n221), .O(n224));
  inv1   g138(.a(n224), .O(n225));
  inv1   g139(.a(G171gat), .O(n226));
  nor2   g140(.a(G177gat), .b(n226), .O(n227));
  inv1   g141(.a(G177gat), .O(n228));
  nor2   g142(.a(n228), .b(G171gat), .O(n229));
  nor2   g143(.a(n229), .b(n227), .O(n230));
  nor2   g144(.a(n230), .b(n181), .O(n231));
  inv1   g145(.a(n230), .O(n232));
  nor2   g146(.a(n232), .b(G130gat), .O(n233));
  nor2   g147(.a(n233), .b(n231), .O(n234));
  nor2   g148(.a(n234), .b(n225), .O(n235));
  inv1   g149(.a(n234), .O(n236));
  nor2   g150(.a(n236), .b(n224), .O(n237));
  nor2   g151(.a(n237), .b(n235), .O(n238));
  inv1   g152(.a(n238), .O(n239));
  nor2   g153(.a(n239), .b(n214), .O(n240));
  nor2   g154(.a(n238), .b(n213), .O(n241));
  nor2   g155(.a(n241), .b(n240), .O(G768gat));
  inv1   g156(.a(G153gat), .O(n243));
  inv1   g157(.a(G447gat), .O(n244));
  inv1   g158(.a(G156gat), .O(n245));
  nor2   g159(.a(n245), .b(n118), .O(n246));
  nor2   g160(.a(n246), .b(n244), .O(n247));
  inv1   g161(.a(n247), .O(n248));
  nor2   g162(.a(n248), .b(n103), .O(n249));
  nor2   g163(.a(n249), .b(n106), .O(n250));
  nor2   g164(.a(n250), .b(n243), .O(n251));
  nor2   g165(.a(n120), .b(n87), .O(n252));
  nor2   g166(.a(n135), .b(n103), .O(n253));
  inv1   g167(.a(n253), .O(n254));
  nor2   g168(.a(n254), .b(n109), .O(n255));
  inv1   g169(.a(n255), .O(n256));
  nor2   g170(.a(n256), .b(n252), .O(n257));
  nor2   g171(.a(G42gat), .b(n103), .O(n258));
  nor2   g172(.a(n87), .b(G17gat), .O(n259));
  nor2   g173(.a(n259), .b(n258), .O(n260));
  inv1   g174(.a(n246), .O(n261));
  nor2   g175(.a(n261), .b(n244), .O(n262));
  inv1   g176(.a(n262), .O(n263));
  nor2   g177(.a(n263), .b(n260), .O(n264));
  nor2   g178(.a(n264), .b(n257), .O(n265));
  nor2   g179(.a(n265), .b(n162), .O(n266));
  nor2   g180(.a(n91), .b(n93), .O(n267));
  inv1   g181(.a(n267), .O(n268));
  nor2   g182(.a(n268), .b(n244), .O(n269));
  inv1   g183(.a(n269), .O(n270));
  nor2   g184(.a(G268gat), .b(n137), .O(n271));
  inv1   g185(.a(n271), .O(n272));
  nor2   g186(.a(n272), .b(n270), .O(n273));
  nor2   g187(.a(n273), .b(n266), .O(n274));
  inv1   g188(.a(n274), .O(n275));
  nor2   g189(.a(n275), .b(n251), .O(n276));
  nor2   g190(.a(n276), .b(n207), .O(n277));
  inv1   g191(.a(G261gat), .O(n278));
  inv1   g192(.a(n276), .O(n279));
  nor2   g193(.a(n279), .b(G201gat), .O(n280));
  nor2   g194(.a(n280), .b(n278), .O(n281));
  inv1   g195(.a(n281), .O(n282));
  nor2   g196(.a(n282), .b(n277), .O(n283));
  inv1   g197(.a(G219gat), .O(n284));
  nor2   g198(.a(n280), .b(n277), .O(n285));
  nor2   g199(.a(n285), .b(G261gat), .O(n286));
  nor2   g200(.a(n286), .b(n284), .O(n287));
  inv1   g201(.a(n287), .O(n288));
  nor2   g202(.a(n288), .b(n283), .O(n289));
  inv1   g203(.a(G228gat), .O(n290));
  inv1   g204(.a(n285), .O(n291));
  nor2   g205(.a(n291), .b(n290), .O(n292));
  inv1   g206(.a(G237gat), .O(n293));
  inv1   g207(.a(n277), .O(n294));
  nor2   g208(.a(n294), .b(n293), .O(n295));
  inv1   g209(.a(G246gat), .O(n296));
  nor2   g210(.a(n276), .b(n296), .O(n297));
  inv1   g211(.a(G73gat), .O(n298));
  inv1   g212(.a(G72gat), .O(n299));
  nor2   g213(.a(n299), .b(n87), .O(n300));
  inv1   g214(.a(n300), .O(n301));
  nor2   g215(.a(n301), .b(n298), .O(n302));
  inv1   g216(.a(n302), .O(n303));
  nor2   g217(.a(n303), .b(n150), .O(n304));
  inv1   g218(.a(n304), .O(n305));
  nor2   g219(.a(n305), .b(n207), .O(n306));
  inv1   g220(.a(G210gat), .O(n307));
  nor2   g221(.a(n307), .b(n160), .O(n308));
  inv1   g222(.a(G255gat), .O(n309));
  inv1   g223(.a(G267gat), .O(n310));
  nor2   g224(.a(n310), .b(n309), .O(n311));
  nor2   g225(.a(n311), .b(n308), .O(n312));
  inv1   g226(.a(n312), .O(n313));
  nor2   g227(.a(n313), .b(n306), .O(n314));
  inv1   g228(.a(n314), .O(n315));
  nor2   g229(.a(n315), .b(n297), .O(n316));
  inv1   g230(.a(n316), .O(n317));
  nor2   g231(.a(n317), .b(n295), .O(n318));
  inv1   g232(.a(n318), .O(n319));
  nor2   g233(.a(n319), .b(n292), .O(n320));
  inv1   g234(.a(n320), .O(n321));
  nor2   g235(.a(n321), .b(n289), .O(n322));
  inv1   g236(.a(n322), .O(G850gat));
  nor2   g237(.a(n265), .b(n171), .O(n324));
  inv1   g238(.a(G143gat), .O(n325));
  nor2   g239(.a(n250), .b(n325), .O(n326));
  nor2   g240(.a(n326), .b(n273), .O(n327));
  inv1   g241(.a(n327), .O(n328));
  nor2   g242(.a(n328), .b(n324), .O(n329));
  inv1   g243(.a(n329), .O(n330));
  nor2   g244(.a(n330), .b(G183gat), .O(n331));
  nor2   g245(.a(n329), .b(n216), .O(n332));
  nor2   g246(.a(n332), .b(n331), .O(n333));
  inv1   g247(.a(n333), .O(n334));
  nor2   g248(.a(n281), .b(n277), .O(n335));
  nor2   g249(.a(n265), .b(n172), .O(n336));
  inv1   g250(.a(G146gat), .O(n337));
  nor2   g251(.a(n250), .b(n337), .O(n338));
  nor2   g252(.a(n338), .b(n273), .O(n339));
  inv1   g253(.a(n339), .O(n340));
  nor2   g254(.a(n340), .b(n336), .O(n341));
  inv1   g255(.a(n341), .O(n342));
  nor2   g256(.a(n342), .b(G189gat), .O(n343));
  nor2   g257(.a(n265), .b(n160), .O(n344));
  inv1   g258(.a(G149gat), .O(n345));
  nor2   g259(.a(n250), .b(n345), .O(n346));
  nor2   g260(.a(n346), .b(n273), .O(n347));
  inv1   g261(.a(n347), .O(n348));
  nor2   g262(.a(n348), .b(n344), .O(n349));
  inv1   g263(.a(n349), .O(n350));
  nor2   g264(.a(n350), .b(G195gat), .O(n351));
  nor2   g265(.a(n351), .b(n343), .O(n352));
  inv1   g266(.a(n352), .O(n353));
  nor2   g267(.a(n353), .b(n335), .O(n354));
  nor2   g268(.a(n341), .b(n217), .O(n355));
  nor2   g269(.a(n349), .b(n205), .O(n356));
  inv1   g270(.a(n356), .O(n357));
  nor2   g271(.a(n357), .b(n343), .O(n358));
  nor2   g272(.a(n358), .b(n355), .O(n359));
  inv1   g273(.a(n359), .O(n360));
  nor2   g274(.a(n360), .b(n354), .O(n361));
  nor2   g275(.a(n361), .b(n334), .O(n362));
  inv1   g276(.a(n361), .O(n363));
  nor2   g277(.a(n363), .b(n333), .O(n364));
  nor2   g278(.a(n364), .b(n284), .O(n365));
  inv1   g279(.a(n365), .O(n366));
  nor2   g280(.a(n366), .b(n362), .O(n367));
  nor2   g281(.a(n334), .b(n290), .O(n368));
  inv1   g282(.a(n332), .O(n369));
  nor2   g283(.a(n369), .b(n293), .O(n370));
  nor2   g284(.a(n329), .b(n296), .O(n371));
  nor2   g285(.a(n305), .b(n216), .O(n372));
  nor2   g286(.a(n307), .b(n184), .O(n373));
  nor2   g287(.a(n373), .b(n372), .O(n374));
  inv1   g288(.a(n374), .O(n375));
  nor2   g289(.a(n375), .b(n371), .O(n376));
  inv1   g290(.a(n376), .O(n377));
  nor2   g291(.a(n377), .b(n370), .O(n378));
  inv1   g292(.a(n378), .O(n379));
  nor2   g293(.a(n379), .b(n368), .O(n380));
  inv1   g294(.a(n380), .O(n381));
  nor2   g295(.a(n381), .b(n367), .O(n382));
  inv1   g296(.a(n382), .O(G863gat));
  nor2   g297(.a(n355), .b(n343), .O(n384));
  nor2   g298(.a(n351), .b(n335), .O(n385));
  nor2   g299(.a(n385), .b(n356), .O(n386));
  inv1   g300(.a(n386), .O(n387));
  nor2   g301(.a(n387), .b(n384), .O(n388));
  inv1   g302(.a(n384), .O(n389));
  nor2   g303(.a(n386), .b(n389), .O(n390));
  nor2   g304(.a(n390), .b(n284), .O(n391));
  inv1   g305(.a(n391), .O(n392));
  nor2   g306(.a(n392), .b(n388), .O(n393));
  nor2   g307(.a(n389), .b(n290), .O(n394));
  inv1   g308(.a(n355), .O(n395));
  nor2   g309(.a(n395), .b(n293), .O(n396));
  nor2   g310(.a(n341), .b(n296), .O(n397));
  nor2   g311(.a(n305), .b(n217), .O(n398));
  nor2   g312(.a(n307), .b(n171), .O(n399));
  inv1   g313(.a(G259gat), .O(n400));
  nor2   g314(.a(n400), .b(n309), .O(n401));
  nor2   g315(.a(n401), .b(n399), .O(n402));
  inv1   g316(.a(n402), .O(n403));
  nor2   g317(.a(n403), .b(n398), .O(n404));
  inv1   g318(.a(n404), .O(n405));
  nor2   g319(.a(n405), .b(n397), .O(n406));
  inv1   g320(.a(n406), .O(n407));
  nor2   g321(.a(n407), .b(n396), .O(n408));
  inv1   g322(.a(n408), .O(n409));
  nor2   g323(.a(n409), .b(n394), .O(n410));
  inv1   g324(.a(n410), .O(n411));
  nor2   g325(.a(n411), .b(n393), .O(n412));
  inv1   g326(.a(n412), .O(G864gat));
  nor2   g327(.a(n356), .b(n351), .O(n414));
  inv1   g328(.a(n414), .O(n415));
  nor2   g329(.a(n415), .b(n335), .O(n416));
  inv1   g330(.a(n335), .O(n417));
  nor2   g331(.a(n414), .b(n417), .O(n418));
  nor2   g332(.a(n418), .b(n284), .O(n419));
  inv1   g333(.a(n419), .O(n420));
  nor2   g334(.a(n420), .b(n416), .O(n421));
  nor2   g335(.a(n415), .b(n290), .O(n422));
  nor2   g336(.a(n357), .b(n293), .O(n423));
  nor2   g337(.a(n349), .b(n296), .O(n424));
  nor2   g338(.a(n305), .b(n205), .O(n425));
  nor2   g339(.a(n307), .b(n172), .O(n426));
  inv1   g340(.a(G260gat), .O(n427));
  nor2   g341(.a(n427), .b(n309), .O(n428));
  nor2   g342(.a(n428), .b(n426), .O(n429));
  inv1   g343(.a(n429), .O(n430));
  nor2   g344(.a(n430), .b(n425), .O(n431));
  inv1   g345(.a(n431), .O(n432));
  nor2   g346(.a(n432), .b(n424), .O(n433));
  inv1   g347(.a(n433), .O(n434));
  nor2   g348(.a(n434), .b(n423), .O(n435));
  inv1   g349(.a(n435), .O(n436));
  nor2   g350(.a(n436), .b(n422), .O(n437));
  inv1   g351(.a(n437), .O(n438));
  nor2   g352(.a(n438), .b(n421), .O(n439));
  inv1   g353(.a(n439), .O(G865gat));
  nor2   g354(.a(n265), .b(n154), .O(n441));
  nor2   g355(.a(n248), .b(n137), .O(n442));
  inv1   g356(.a(n442), .O(n443));
  nor2   g357(.a(n443), .b(n325), .O(n444));
  inv1   g358(.a(G138gat), .O(n445));
  nor2   g359(.a(n445), .b(n107), .O(n446));
  nor2   g360(.a(G268gat), .b(n103), .O(n447));
  inv1   g361(.a(n447), .O(n448));
  nor2   g362(.a(n448), .b(n270), .O(n449));
  nor2   g363(.a(n449), .b(n446), .O(n450));
  inv1   g364(.a(n450), .O(n451));
  nor2   g365(.a(n451), .b(n444), .O(n452));
  inv1   g366(.a(n452), .O(n453));
  nor2   g367(.a(n453), .b(n441), .O(n454));
  nor2   g368(.a(n454), .b(n199), .O(n455));
  inv1   g369(.a(n454), .O(n456));
  nor2   g370(.a(n456), .b(G159gat), .O(n457));
  nor2   g371(.a(n265), .b(n184), .O(n458));
  nor2   g372(.a(n443), .b(n243), .O(n459));
  inv1   g373(.a(G152gat), .O(n460));
  nor2   g374(.a(n460), .b(n445), .O(n461));
  nor2   g375(.a(n461), .b(n449), .O(n462));
  inv1   g376(.a(n462), .O(n463));
  nor2   g377(.a(n463), .b(n459), .O(n464));
  inv1   g378(.a(n464), .O(n465));
  nor2   g379(.a(n465), .b(n458), .O(n466));
  inv1   g380(.a(n466), .O(n467));
  nor2   g381(.a(n467), .b(G177gat), .O(n468));
  nor2   g382(.a(n361), .b(n331), .O(n469));
  nor2   g383(.a(n469), .b(n332), .O(n470));
  nor2   g384(.a(n470), .b(n468), .O(n471));
  inv1   g385(.a(n471), .O(n472));
  nor2   g386(.a(n265), .b(n155), .O(n473));
  nor2   g387(.a(n443), .b(n337), .O(n474));
  nor2   g388(.a(n445), .b(n135), .O(n475));
  nor2   g389(.a(n475), .b(n449), .O(n476));
  inv1   g390(.a(n476), .O(n477));
  nor2   g391(.a(n477), .b(n474), .O(n478));
  inv1   g392(.a(n478), .O(n479));
  nor2   g393(.a(n479), .b(n473), .O(n480));
  inv1   g394(.a(n480), .O(n481));
  nor2   g395(.a(n481), .b(G165gat), .O(n482));
  nor2   g396(.a(n265), .b(n182), .O(n483));
  nor2   g397(.a(n443), .b(n345), .O(n484));
  nor2   g398(.a(n445), .b(n103), .O(n485));
  nor2   g399(.a(n485), .b(n449), .O(n486));
  inv1   g400(.a(n486), .O(n487));
  nor2   g401(.a(n487), .b(n484), .O(n488));
  inv1   g402(.a(n488), .O(n489));
  nor2   g403(.a(n489), .b(n483), .O(n490));
  inv1   g404(.a(n490), .O(n491));
  nor2   g405(.a(n491), .b(G171gat), .O(n492));
  nor2   g406(.a(n492), .b(n482), .O(n493));
  inv1   g407(.a(n493), .O(n494));
  nor2   g408(.a(n494), .b(n472), .O(n495));
  nor2   g409(.a(n480), .b(n200), .O(n496));
  nor2   g410(.a(n466), .b(n228), .O(n497));
  nor2   g411(.a(n490), .b(n226), .O(n498));
  nor2   g412(.a(n498), .b(n497), .O(n499));
  nor2   g413(.a(n499), .b(n492), .O(n500));
  inv1   g414(.a(n500), .O(n501));
  nor2   g415(.a(n501), .b(n482), .O(n502));
  nor2   g416(.a(n502), .b(n496), .O(n503));
  inv1   g417(.a(n503), .O(n504));
  nor2   g418(.a(n504), .b(n495), .O(n505));
  nor2   g419(.a(n505), .b(n457), .O(n506));
  nor2   g420(.a(n506), .b(n455), .O(n507));
  inv1   g421(.a(n507), .O(G866gat));
  nor2   g422(.a(n497), .b(n468), .O(n509));
  inv1   g423(.a(n509), .O(n510));
  nor2   g424(.a(n510), .b(n470), .O(n511));
  inv1   g425(.a(n470), .O(n512));
  nor2   g426(.a(n509), .b(n512), .O(n513));
  nor2   g427(.a(n513), .b(n284), .O(n514));
  inv1   g428(.a(n514), .O(n515));
  nor2   g429(.a(n515), .b(n511), .O(n516));
  nor2   g430(.a(n510), .b(n290), .O(n517));
  inv1   g431(.a(n497), .O(n518));
  nor2   g432(.a(n518), .b(n293), .O(n519));
  nor2   g433(.a(n466), .b(n296), .O(n520));
  nor2   g434(.a(n305), .b(n228), .O(n521));
  nor2   g435(.a(n307), .b(n182), .O(n522));
  nor2   g436(.a(n522), .b(n521), .O(n523));
  inv1   g437(.a(n523), .O(n524));
  nor2   g438(.a(n524), .b(n520), .O(n525));
  inv1   g439(.a(n525), .O(n526));
  nor2   g440(.a(n526), .b(n519), .O(n527));
  inv1   g441(.a(n527), .O(n528));
  nor2   g442(.a(n528), .b(n517), .O(n529));
  inv1   g443(.a(n529), .O(n530));
  nor2   g444(.a(n530), .b(n516), .O(n531));
  inv1   g445(.a(n531), .O(G874gat));
  nor2   g446(.a(n457), .b(n455), .O(n533));
  inv1   g447(.a(n533), .O(n534));
  nor2   g448(.a(n534), .b(n505), .O(n535));
  inv1   g449(.a(n505), .O(n536));
  nor2   g450(.a(n533), .b(n536), .O(n537));
  nor2   g451(.a(n537), .b(n284), .O(n538));
  inv1   g452(.a(n538), .O(n539));
  nor2   g453(.a(n539), .b(n535), .O(n540));
  nor2   g454(.a(n534), .b(n290), .O(n541));
  inv1   g455(.a(n455), .O(n542));
  nor2   g456(.a(n542), .b(n293), .O(n543));
  nor2   g457(.a(n454), .b(n296), .O(n544));
  nor2   g458(.a(n305), .b(n199), .O(n545));
  inv1   g459(.a(G268gat), .O(n546));
  nor2   g460(.a(n546), .b(n307), .O(n547));
  nor2   g461(.a(n547), .b(n545), .O(n548));
  inv1   g462(.a(n548), .O(n549));
  nor2   g463(.a(n549), .b(n544), .O(n550));
  inv1   g464(.a(n550), .O(n551));
  nor2   g465(.a(n551), .b(n543), .O(n552));
  inv1   g466(.a(n552), .O(n553));
  nor2   g467(.a(n553), .b(n541), .O(n554));
  inv1   g468(.a(n554), .O(n555));
  nor2   g469(.a(n555), .b(n540), .O(n556));
  inv1   g470(.a(n556), .O(G878gat));
  nor2   g471(.a(n496), .b(n482), .O(n558));
  nor2   g472(.a(n492), .b(n472), .O(n559));
  nor2   g473(.a(n559), .b(n500), .O(n560));
  inv1   g474(.a(n560), .O(n561));
  nor2   g475(.a(n561), .b(n558), .O(n562));
  inv1   g476(.a(n558), .O(n563));
  nor2   g477(.a(n560), .b(n563), .O(n564));
  nor2   g478(.a(n564), .b(n284), .O(n565));
  inv1   g479(.a(n565), .O(n566));
  nor2   g480(.a(n566), .b(n562), .O(n567));
  nor2   g481(.a(n563), .b(n290), .O(n568));
  inv1   g482(.a(n496), .O(n569));
  nor2   g483(.a(n569), .b(n293), .O(n570));
  nor2   g484(.a(n480), .b(n296), .O(n571));
  nor2   g485(.a(n305), .b(n200), .O(n572));
  nor2   g486(.a(n307), .b(n154), .O(n573));
  nor2   g487(.a(n573), .b(n572), .O(n574));
  inv1   g488(.a(n574), .O(n575));
  nor2   g489(.a(n575), .b(n571), .O(n576));
  inv1   g490(.a(n576), .O(n577));
  nor2   g491(.a(n577), .b(n570), .O(n578));
  inv1   g492(.a(n578), .O(n579));
  nor2   g493(.a(n579), .b(n568), .O(n580));
  inv1   g494(.a(n580), .O(n581));
  nor2   g495(.a(n581), .b(n567), .O(n582));
  inv1   g496(.a(n582), .O(G879gat));
  nor2   g497(.a(n498), .b(n492), .O(n584));
  nor2   g498(.a(n497), .b(n471), .O(n585));
  inv1   g499(.a(n585), .O(n586));
  nor2   g500(.a(n586), .b(n584), .O(n587));
  inv1   g501(.a(n584), .O(n588));
  nor2   g502(.a(n585), .b(n588), .O(n589));
  nor2   g503(.a(n589), .b(n284), .O(n590));
  inv1   g504(.a(n590), .O(n591));
  nor2   g505(.a(n591), .b(n587), .O(n592));
  nor2   g506(.a(n588), .b(n290), .O(n593));
  inv1   g507(.a(n498), .O(n594));
  nor2   g508(.a(n594), .b(n293), .O(n595));
  nor2   g509(.a(n490), .b(n296), .O(n596));
  nor2   g510(.a(n305), .b(n226), .O(n597));
  nor2   g511(.a(n307), .b(n155), .O(n598));
  nor2   g512(.a(n598), .b(n597), .O(n599));
  inv1   g513(.a(n599), .O(n600));
  nor2   g514(.a(n600), .b(n596), .O(n601));
  inv1   g515(.a(n601), .O(n602));
  nor2   g516(.a(n602), .b(n595), .O(n603));
  inv1   g517(.a(n603), .O(n604));
  nor2   g518(.a(n604), .b(n593), .O(n605));
  inv1   g519(.a(n605), .O(n606));
  nor2   g520(.a(n606), .b(n592), .O(n607));
  inv1   g521(.a(n607), .O(G880gat));
endmodule


