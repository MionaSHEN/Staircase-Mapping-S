// Benchmark "c3540_blif" written by ABC on Sun Apr 14 20:12:58 2019

module c3540_blif  ( 
    G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
    G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200,
    G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274,
    G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698,
    G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107,
    G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
    G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270,
    G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire n73, n74, n75, n76, n78, n79, n80, n82, n83, n84, n85, n86, n87, n88,
    n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n142, n143, n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
    n163, n164, n165, n166, n167, n168, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n194, n195, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
    n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
    n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n790, n791, n792, n793,
    n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
    n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n870, n871, n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
    n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
    n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
    n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
    n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
    n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
    n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
    n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
    n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1190, n1191, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
    n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
    n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
    n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
    n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
    n1273, n1274, n1275, n1276, n1277, n1278, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
    n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
    n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
    n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
    n1425, n1426, n1427, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1452, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1483, n1484;
  nor2   g0000(.a(G58), .b(G50), .O(n73));
  inv1   g0001(.a(n73), .O(n74));
  nor2   g0002(.a(n74), .b(G68), .O(n75));
  inv1   g0003(.a(n75), .O(n76));
  nor2   g0004(.a(n76), .b(G77), .O(G353));
  inv1   g0005(.a(G87), .O(n78));
  nor2   g0006(.a(G107), .b(G97), .O(n79));
  nor2   g0007(.a(n79), .b(n78), .O(n80));
  inv1   g0008(.a(n80), .O(G355));
  inv1   g0009(.a(G1), .O(n82));
  inv1   g0010(.a(G20), .O(n83));
  nor2   g0011(.a(n83), .b(n82), .O(n84));
  inv1   g0012(.a(G77), .O(n85));
  inv1   g0013(.a(G244), .O(n86));
  nor2   g0014(.a(n86), .b(n85), .O(n87));
  inv1   g0015(.a(G116), .O(n88));
  inv1   g0016(.a(G270), .O(n89));
  nor2   g0017(.a(n89), .b(n88), .O(n90));
  nor2   g0018(.a(n90), .b(n87), .O(n91));
  inv1   g0019(.a(n91), .O(n92));
  inv1   g0020(.a(G58), .O(n93));
  inv1   g0021(.a(G232), .O(n94));
  nor2   g0022(.a(n94), .b(n93), .O(n95));
  inv1   g0023(.a(G97), .O(n96));
  inv1   g0024(.a(G257), .O(n97));
  nor2   g0025(.a(n97), .b(n96), .O(n98));
  nor2   g0026(.a(n98), .b(n95), .O(n99));
  inv1   g0027(.a(n99), .O(n100));
  nor2   g0028(.a(n100), .b(n92), .O(n101));
  inv1   g0029(.a(n101), .O(n102));
  inv1   g0030(.a(G107), .O(n103));
  inv1   g0031(.a(G264), .O(n104));
  nor2   g0032(.a(n104), .b(n103), .O(n105));
  inv1   g0033(.a(G50), .O(n106));
  inv1   g0034(.a(G226), .O(n107));
  nor2   g0035(.a(n107), .b(n106), .O(n108));
  nor2   g0036(.a(n108), .b(n105), .O(n109));
  inv1   g0037(.a(n109), .O(n110));
  inv1   g0038(.a(G68), .O(n111));
  inv1   g0039(.a(G238), .O(n112));
  nor2   g0040(.a(n112), .b(n111), .O(n113));
  inv1   g0041(.a(G250), .O(n114));
  nor2   g0042(.a(n114), .b(n78), .O(n115));
  nor2   g0043(.a(n115), .b(n113), .O(n116));
  inv1   g0044(.a(n116), .O(n117));
  nor2   g0045(.a(n117), .b(n110), .O(n118));
  inv1   g0046(.a(n118), .O(n119));
  nor2   g0047(.a(n119), .b(n102), .O(n120));
  nor2   g0048(.a(n120), .b(n84), .O(n121));
  inv1   g0049(.a(G13), .O(n122));
  nor2   g0050(.a(n122), .b(n82), .O(n123));
  inv1   g0051(.a(n123), .O(n124));
  nor2   g0052(.a(n124), .b(n83), .O(n125));
  inv1   g0053(.a(n125), .O(n126));
  nor2   g0054(.a(G68), .b(G58), .O(n127));
  nor2   g0055(.a(n127), .b(n106), .O(n128));
  inv1   g0056(.a(n128), .O(n129));
  nor2   g0057(.a(n129), .b(n126), .O(n130));
  nor2   g0058(.a(G13), .b(n82), .O(n131));
  inv1   g0059(.a(n131), .O(n132));
  nor2   g0060(.a(n132), .b(n83), .O(n133));
  inv1   g0061(.a(n133), .O(n134));
  nor2   g0062(.a(G264), .b(G257), .O(n135));
  nor2   g0063(.a(n135), .b(n114), .O(n136));
  inv1   g0064(.a(n136), .O(n137));
  nor2   g0065(.a(n137), .b(n134), .O(n138));
  nor2   g0066(.a(n138), .b(n130), .O(n139));
  inv1   g0067(.a(n139), .O(n140));
  nor2   g0068(.a(n140), .b(n121), .O(G361));
  nor2   g0069(.a(n89), .b(G264), .O(n142));
  nor2   g0070(.a(G270), .b(n104), .O(n143));
  nor2   g0071(.a(n143), .b(n142), .O(n144));
  nor2   g0072(.a(n144), .b(n114), .O(n145));
  inv1   g0073(.a(n144), .O(n146));
  nor2   g0074(.a(n146), .b(G250), .O(n147));
  nor2   g0075(.a(n147), .b(n145), .O(n148));
  inv1   g0076(.a(n148), .O(n149));
  nor2   g0077(.a(n149), .b(n97), .O(n150));
  nor2   g0078(.a(n148), .b(G257), .O(n151));
  nor2   g0079(.a(n151), .b(n150), .O(n152));
  inv1   g0080(.a(n152), .O(n153));
  nor2   g0081(.a(n86), .b(G238), .O(n154));
  nor2   g0082(.a(G244), .b(n112), .O(n155));
  nor2   g0083(.a(n155), .b(n154), .O(n156));
  nor2   g0084(.a(n156), .b(n107), .O(n157));
  inv1   g0085(.a(n156), .O(n158));
  nor2   g0086(.a(n158), .b(G226), .O(n159));
  nor2   g0087(.a(n159), .b(n157), .O(n160));
  inv1   g0088(.a(n160), .O(n161));
  nor2   g0089(.a(n161), .b(n94), .O(n162));
  nor2   g0090(.a(n160), .b(G232), .O(n163));
  nor2   g0091(.a(n163), .b(n162), .O(n164));
  inv1   g0092(.a(n164), .O(n165));
  nor2   g0093(.a(n165), .b(n153), .O(n166));
  nor2   g0094(.a(n164), .b(n152), .O(n167));
  nor2   g0095(.a(n167), .b(n166), .O(n168));
  inv1   g0096(.a(n168), .O(G358));
  nor2   g0097(.a(n103), .b(G97), .O(n170));
  nor2   g0098(.a(G107), .b(n96), .O(n171));
  nor2   g0099(.a(n171), .b(n170), .O(n172));
  nor2   g0100(.a(G116), .b(n78), .O(n173));
  nor2   g0101(.a(n88), .b(G87), .O(n174));
  nor2   g0102(.a(n174), .b(n173), .O(n175));
  inv1   g0103(.a(n175), .O(n176));
  nor2   g0104(.a(n176), .b(n172), .O(n177));
  inv1   g0105(.a(n172), .O(n178));
  nor2   g0106(.a(n175), .b(n178), .O(n179));
  nor2   g0107(.a(n179), .b(n177), .O(n180));
  inv1   g0108(.a(n180), .O(n181));
  nor2   g0109(.a(n111), .b(G58), .O(n182));
  nor2   g0110(.a(G68), .b(n93), .O(n183));
  nor2   g0111(.a(n183), .b(n182), .O(n184));
  nor2   g0112(.a(n184), .b(n85), .O(n185));
  inv1   g0113(.a(n184), .O(n186));
  nor2   g0114(.a(n186), .b(G77), .O(n187));
  nor2   g0115(.a(n187), .b(n185), .O(n188));
  inv1   g0116(.a(n188), .O(n189));
  nor2   g0117(.a(n189), .b(n106), .O(n190));
  nor2   g0118(.a(n188), .b(G50), .O(n191));
  nor2   g0119(.a(n191), .b(n190), .O(n192));
  inv1   g0120(.a(n192), .O(n193));
  nor2   g0121(.a(n193), .b(n181), .O(n194));
  nor2   g0122(.a(n192), .b(n180), .O(n195));
  nor2   g0123(.a(n195), .b(n194), .O(G351));
  inv1   g0124(.a(G33), .O(n197));
  inv1   g0125(.a(G41), .O(n198));
  nor2   g0126(.a(n198), .b(n197), .O(n199));
  nor2   g0127(.a(n199), .b(n124), .O(n200));
  inv1   g0128(.a(n200), .O(n201));
  nor2   g0129(.a(G1698), .b(G33), .O(n202));
  nor2   g0130(.a(n202), .b(G33), .O(n203));
  inv1   g0131(.a(n203), .O(n204));
  nor2   g0132(.a(n204), .b(n86), .O(n205));
  nor2   g0133(.a(n88), .b(n197), .O(n206));
  inv1   g0134(.a(n202), .O(n207));
  nor2   g0135(.a(n207), .b(n112), .O(n208));
  nor2   g0136(.a(n208), .b(n206), .O(n209));
  inv1   g0137(.a(n209), .O(n210));
  nor2   g0138(.a(n210), .b(n205), .O(n211));
  nor2   g0139(.a(n211), .b(n201), .O(n212));
  inv1   g0140(.a(G274), .O(n213));
  nor2   g0141(.a(n200), .b(n213), .O(n214));
  inv1   g0142(.a(n214), .O(n215));
  inv1   g0143(.a(G45), .O(n216));
  nor2   g0144(.a(n216), .b(G1), .O(n217));
  inv1   g0145(.a(n217), .O(n218));
  nor2   g0146(.a(n218), .b(n215), .O(n219));
  nor2   g0147(.a(n217), .b(n114), .O(n220));
  inv1   g0148(.a(n220), .O(n221));
  nor2   g0149(.a(n221), .b(n200), .O(n222));
  nor2   g0150(.a(n222), .b(n219), .O(n223));
  inv1   g0151(.a(n223), .O(n224));
  nor2   g0152(.a(n224), .b(n212), .O(n225));
  inv1   g0153(.a(n225), .O(n226));
  nor2   g0154(.a(n226), .b(G179), .O(n227));
  nor2   g0155(.a(n225), .b(G169), .O(n228));
  inv1   g0156(.a(n84), .O(n229));
  nor2   g0157(.a(n229), .b(n197), .O(n230));
  nor2   g0158(.a(n230), .b(n123), .O(n231));
  nor2   g0159(.a(G33), .b(G20), .O(n232));
  inv1   g0160(.a(n232), .O(n233));
  nor2   g0161(.a(n233), .b(n111), .O(n234));
  nor2   g0162(.a(n197), .b(G20), .O(n235));
  inv1   g0163(.a(n235), .O(n236));
  nor2   g0164(.a(n236), .b(n96), .O(n237));
  nor2   g0165(.a(G97), .b(G87), .O(n238));
  inv1   g0166(.a(n238), .O(n239));
  nor2   g0167(.a(n239), .b(G107), .O(n240));
  nor2   g0168(.a(n240), .b(n83), .O(n241));
  nor2   g0169(.a(n241), .b(n237), .O(n242));
  inv1   g0170(.a(n242), .O(n243));
  nor2   g0171(.a(n243), .b(n234), .O(n244));
  nor2   g0172(.a(n244), .b(n231), .O(n245));
  nor2   g0173(.a(n122), .b(G1), .O(n246));
  inv1   g0174(.a(n246), .O(n247));
  nor2   g0175(.a(n247), .b(n83), .O(n248));
  nor2   g0176(.a(n197), .b(G1), .O(n249));
  nor2   g0177(.a(n249), .b(n78), .O(n250));
  nor2   g0178(.a(n250), .b(n248), .O(n251));
  inv1   g0179(.a(n231), .O(n252));
  nor2   g0180(.a(n248), .b(n252), .O(n253));
  nor2   g0181(.a(n253), .b(n78), .O(n254));
  nor2   g0182(.a(n254), .b(n251), .O(n255));
  nor2   g0183(.a(n255), .b(n245), .O(n256));
  nor2   g0184(.a(n256), .b(n228), .O(n257));
  inv1   g0185(.a(n257), .O(n258));
  nor2   g0186(.a(n258), .b(n227), .O(n259));
  inv1   g0187(.a(G200), .O(n260));
  nor2   g0188(.a(n225), .b(n260), .O(n261));
  inv1   g0189(.a(n256), .O(n262));
  inv1   g0190(.a(G190), .O(n263));
  nor2   g0191(.a(n226), .b(n263), .O(n264));
  nor2   g0192(.a(n264), .b(n262), .O(n265));
  inv1   g0193(.a(n265), .O(n266));
  nor2   g0194(.a(n266), .b(n261), .O(n267));
  nor2   g0195(.a(n267), .b(n259), .O(n268));
  inv1   g0196(.a(n268), .O(n269));
  nor2   g0197(.a(n204), .b(n114), .O(n270));
  nor2   g0198(.a(n207), .b(n86), .O(n271));
  inv1   g0199(.a(G283), .O(n272));
  nor2   g0200(.a(n272), .b(n197), .O(n273));
  nor2   g0201(.a(n273), .b(n271), .O(n274));
  inv1   g0202(.a(n274), .O(n275));
  nor2   g0203(.a(n275), .b(n270), .O(n276));
  nor2   g0204(.a(n276), .b(n201), .O(n277));
  nor2   g0205(.a(n218), .b(G41), .O(n278));
  inv1   g0206(.a(n278), .O(n279));
  nor2   g0207(.a(n279), .b(n215), .O(n280));
  nor2   g0208(.a(n278), .b(n200), .O(n281));
  inv1   g0209(.a(n281), .O(n282));
  nor2   g0210(.a(n282), .b(n97), .O(n283));
  nor2   g0211(.a(n283), .b(n280), .O(n284));
  inv1   g0212(.a(n284), .O(n285));
  nor2   g0213(.a(n285), .b(n277), .O(n286));
  inv1   g0214(.a(n286), .O(n287));
  nor2   g0215(.a(n287), .b(G179), .O(n288));
  nor2   g0216(.a(n286), .b(G169), .O(n289));
  nor2   g0217(.a(n178), .b(n83), .O(n290));
  nor2   g0218(.a(n233), .b(n85), .O(n291));
  nor2   g0219(.a(n103), .b(n197), .O(n292));
  inv1   g0220(.a(n292), .O(n293));
  nor2   g0221(.a(n293), .b(G20), .O(n294));
  nor2   g0222(.a(n294), .b(n291), .O(n295));
  inv1   g0223(.a(n295), .O(n296));
  nor2   g0224(.a(n296), .b(n290), .O(n297));
  nor2   g0225(.a(n297), .b(n231), .O(n298));
  nor2   g0226(.a(n249), .b(n96), .O(n299));
  nor2   g0227(.a(n299), .b(n248), .O(n300));
  nor2   g0228(.a(n253), .b(n96), .O(n301));
  nor2   g0229(.a(n301), .b(n300), .O(n302));
  nor2   g0230(.a(n302), .b(n298), .O(n303));
  nor2   g0231(.a(n303), .b(n289), .O(n304));
  inv1   g0232(.a(n304), .O(n305));
  nor2   g0233(.a(n305), .b(n288), .O(n306));
  nor2   g0234(.a(n286), .b(n260), .O(n307));
  inv1   g0235(.a(n303), .O(n308));
  nor2   g0236(.a(n287), .b(n263), .O(n309));
  nor2   g0237(.a(n309), .b(n308), .O(n310));
  inv1   g0238(.a(n310), .O(n311));
  nor2   g0239(.a(n311), .b(n307), .O(n312));
  nor2   g0240(.a(n312), .b(n306), .O(n313));
  inv1   g0241(.a(n313), .O(n314));
  nor2   g0242(.a(n314), .b(n269), .O(n315));
  inv1   g0243(.a(n315), .O(n316));
  inv1   g0244(.a(G169), .O(n317));
  nor2   g0245(.a(n204), .b(n104), .O(n318));
  nor2   g0246(.a(n207), .b(n97), .O(n319));
  inv1   g0247(.a(G303), .O(n320));
  nor2   g0248(.a(n320), .b(n197), .O(n321));
  nor2   g0249(.a(n321), .b(n319), .O(n322));
  inv1   g0250(.a(n322), .O(n323));
  nor2   g0251(.a(n323), .b(n318), .O(n324));
  nor2   g0252(.a(n324), .b(n201), .O(n325));
  nor2   g0253(.a(n282), .b(n89), .O(n326));
  nor2   g0254(.a(n326), .b(n280), .O(n327));
  inv1   g0255(.a(n327), .O(n328));
  nor2   g0256(.a(n328), .b(n325), .O(n329));
  nor2   g0257(.a(n329), .b(n317), .O(n330));
  inv1   g0258(.a(G179), .O(n331));
  inv1   g0259(.a(n329), .O(n332));
  nor2   g0260(.a(n332), .b(n331), .O(n333));
  nor2   g0261(.a(n333), .b(n330), .O(n334));
  inv1   g0262(.a(n253), .O(n335));
  nor2   g0263(.a(n249), .b(n88), .O(n336));
  inv1   g0264(.a(n336), .O(n337));
  nor2   g0265(.a(n337), .b(n335), .O(n338));
  inv1   g0266(.a(n248), .O(n339));
  nor2   g0267(.a(n339), .b(G116), .O(n340));
  nor2   g0268(.a(n233), .b(n96), .O(n341));
  nor2   g0269(.a(n236), .b(n272), .O(n342));
  nor2   g0270(.a(n88), .b(n83), .O(n343));
  nor2   g0271(.a(n343), .b(n342), .O(n344));
  inv1   g0272(.a(n344), .O(n345));
  nor2   g0273(.a(n345), .b(n341), .O(n346));
  nor2   g0274(.a(n346), .b(n231), .O(n347));
  nor2   g0275(.a(n347), .b(n340), .O(n348));
  inv1   g0276(.a(n348), .O(n349));
  nor2   g0277(.a(n349), .b(n338), .O(n350));
  nor2   g0278(.a(n350), .b(n334), .O(n351));
  nor2   g0279(.a(n329), .b(n260), .O(n352));
  inv1   g0280(.a(n350), .O(n353));
  nor2   g0281(.a(n332), .b(n263), .O(n354));
  nor2   g0282(.a(n354), .b(n353), .O(n355));
  inv1   g0283(.a(n355), .O(n356));
  nor2   g0284(.a(n356), .b(n352), .O(n357));
  nor2   g0285(.a(n357), .b(n351), .O(n358));
  inv1   g0286(.a(n358), .O(n359));
  nor2   g0287(.a(n249), .b(n103), .O(n360));
  inv1   g0288(.a(n360), .O(n361));
  nor2   g0289(.a(n361), .b(n335), .O(n362));
  nor2   g0290(.a(n233), .b(n78), .O(n363));
  nor2   g0291(.a(G107), .b(n83), .O(n364));
  nor2   g0292(.a(n236), .b(n88), .O(n365));
  nor2   g0293(.a(n365), .b(n364), .O(n366));
  inv1   g0294(.a(n366), .O(n367));
  nor2   g0295(.a(n367), .b(n363), .O(n368));
  nor2   g0296(.a(n368), .b(n231), .O(n369));
  nor2   g0297(.a(n339), .b(G107), .O(n370));
  nor2   g0298(.a(n370), .b(n369), .O(n371));
  inv1   g0299(.a(n371), .O(n372));
  nor2   g0300(.a(n372), .b(n362), .O(n373));
  nor2   g0301(.a(n204), .b(n97), .O(n374));
  inv1   g0302(.a(G294), .O(n375));
  nor2   g0303(.a(n375), .b(n197), .O(n376));
  nor2   g0304(.a(n207), .b(n114), .O(n377));
  nor2   g0305(.a(n377), .b(n376), .O(n378));
  inv1   g0306(.a(n378), .O(n379));
  nor2   g0307(.a(n379), .b(n374), .O(n380));
  nor2   g0308(.a(n380), .b(n201), .O(n381));
  nor2   g0309(.a(n282), .b(n104), .O(n382));
  nor2   g0310(.a(n382), .b(n280), .O(n383));
  inv1   g0311(.a(n383), .O(n384));
  nor2   g0312(.a(n384), .b(n381), .O(n385));
  nor2   g0313(.a(n385), .b(G169), .O(n386));
  inv1   g0314(.a(n385), .O(n387));
  nor2   g0315(.a(n387), .b(G179), .O(n388));
  nor2   g0316(.a(n388), .b(n386), .O(n389));
  inv1   g0317(.a(n389), .O(n390));
  nor2   g0318(.a(n390), .b(n373), .O(n391));
  nor2   g0319(.a(n385), .b(n260), .O(n392));
  inv1   g0320(.a(n373), .O(n393));
  nor2   g0321(.a(n387), .b(n263), .O(n394));
  nor2   g0322(.a(n394), .b(n393), .O(n395));
  inv1   g0323(.a(n395), .O(n396));
  nor2   g0324(.a(n396), .b(n392), .O(n397));
  nor2   g0325(.a(n397), .b(n391), .O(n398));
  inv1   g0326(.a(n398), .O(n399));
  nor2   g0327(.a(n399), .b(n359), .O(n400));
  inv1   g0328(.a(n400), .O(n401));
  nor2   g0329(.a(n401), .b(n316), .O(n402));
  inv1   g0330(.a(n402), .O(n403));
  inv1   g0331(.a(G150), .O(n404));
  nor2   g0332(.a(n233), .b(n404), .O(n405));
  nor2   g0333(.a(n75), .b(n83), .O(n406));
  nor2   g0334(.a(n236), .b(n93), .O(n407));
  nor2   g0335(.a(n407), .b(n406), .O(n408));
  inv1   g0336(.a(n408), .O(n409));
  nor2   g0337(.a(n409), .b(n405), .O(n410));
  nor2   g0338(.a(n410), .b(n231), .O(n411));
  nor2   g0339(.a(n339), .b(G50), .O(n412));
  nor2   g0340(.a(n83), .b(G1), .O(n413));
  nor2   g0341(.a(n413), .b(n106), .O(n414));
  inv1   g0342(.a(n414), .O(n415));
  nor2   g0343(.a(n415), .b(n335), .O(n416));
  nor2   g0344(.a(n416), .b(n412), .O(n417));
  inv1   g0345(.a(n417), .O(n418));
  nor2   g0346(.a(n418), .b(n411), .O(n419));
  inv1   g0347(.a(G223), .O(n420));
  nor2   g0348(.a(n204), .b(n420), .O(n421));
  nor2   g0349(.a(n85), .b(n197), .O(n422));
  inv1   g0350(.a(G222), .O(n423));
  nor2   g0351(.a(n207), .b(n423), .O(n424));
  nor2   g0352(.a(n424), .b(n422), .O(n425));
  inv1   g0353(.a(n425), .O(n426));
  nor2   g0354(.a(n426), .b(n421), .O(n427));
  nor2   g0355(.a(n427), .b(n201), .O(n428));
  nor2   g0356(.a(G45), .b(G41), .O(n429));
  nor2   g0357(.a(n429), .b(G1), .O(n430));
  inv1   g0358(.a(n430), .O(n431));
  nor2   g0359(.a(n431), .b(n215), .O(n432));
  nor2   g0360(.a(n430), .b(n200), .O(n433));
  inv1   g0361(.a(n433), .O(n434));
  nor2   g0362(.a(n434), .b(n107), .O(n435));
  nor2   g0363(.a(n435), .b(n432), .O(n436));
  inv1   g0364(.a(n436), .O(n437));
  nor2   g0365(.a(n437), .b(n428), .O(n438));
  nor2   g0366(.a(n438), .b(G169), .O(n439));
  inv1   g0367(.a(n438), .O(n440));
  nor2   g0368(.a(n440), .b(G179), .O(n441));
  nor2   g0369(.a(n441), .b(n439), .O(n442));
  inv1   g0370(.a(n442), .O(n443));
  nor2   g0371(.a(n443), .b(n419), .O(n444));
  nor2   g0372(.a(n438), .b(n260), .O(n445));
  inv1   g0373(.a(n419), .O(n446));
  nor2   g0374(.a(n440), .b(n263), .O(n447));
  nor2   g0375(.a(n447), .b(n446), .O(n448));
  inv1   g0376(.a(n448), .O(n449));
  nor2   g0377(.a(n449), .b(n445), .O(n450));
  nor2   g0378(.a(n450), .b(n444), .O(n451));
  inv1   g0379(.a(n451), .O(n452));
  inv1   g0380(.a(G159), .O(n453));
  nor2   g0381(.a(n233), .b(n453), .O(n454));
  nor2   g0382(.a(n186), .b(n83), .O(n455));
  nor2   g0383(.a(n236), .b(n111), .O(n456));
  nor2   g0384(.a(n456), .b(n455), .O(n457));
  inv1   g0385(.a(n457), .O(n458));
  nor2   g0386(.a(n458), .b(n454), .O(n459));
  nor2   g0387(.a(n459), .b(n231), .O(n460));
  nor2   g0388(.a(n339), .b(G58), .O(n461));
  nor2   g0389(.a(n413), .b(n93), .O(n462));
  inv1   g0390(.a(n462), .O(n463));
  nor2   g0391(.a(n463), .b(n335), .O(n464));
  nor2   g0392(.a(n464), .b(n461), .O(n465));
  inv1   g0393(.a(n465), .O(n466));
  nor2   g0394(.a(n466), .b(n460), .O(n467));
  nor2   g0395(.a(n204), .b(n107), .O(n468));
  nor2   g0396(.a(n207), .b(n420), .O(n469));
  nor2   g0397(.a(n78), .b(n197), .O(n470));
  nor2   g0398(.a(n470), .b(n469), .O(n471));
  inv1   g0399(.a(n471), .O(n472));
  nor2   g0400(.a(n472), .b(n468), .O(n473));
  nor2   g0401(.a(n473), .b(n201), .O(n474));
  nor2   g0402(.a(n434), .b(n94), .O(n475));
  nor2   g0403(.a(n475), .b(n432), .O(n476));
  inv1   g0404(.a(n476), .O(n477));
  nor2   g0405(.a(n477), .b(n474), .O(n478));
  nor2   g0406(.a(n478), .b(G169), .O(n479));
  inv1   g0407(.a(n478), .O(n480));
  nor2   g0408(.a(n480), .b(G179), .O(n481));
  nor2   g0409(.a(n481), .b(n479), .O(n482));
  inv1   g0410(.a(n482), .O(n483));
  nor2   g0411(.a(n483), .b(n467), .O(n484));
  nor2   g0412(.a(n478), .b(n260), .O(n485));
  inv1   g0413(.a(n467), .O(n486));
  nor2   g0414(.a(n480), .b(n263), .O(n487));
  nor2   g0415(.a(n487), .b(n486), .O(n488));
  inv1   g0416(.a(n488), .O(n489));
  nor2   g0417(.a(n489), .b(n485), .O(n490));
  nor2   g0418(.a(n490), .b(n484), .O(n491));
  inv1   g0419(.a(n491), .O(n492));
  nor2   g0420(.a(n492), .b(n452), .O(n493));
  inv1   g0421(.a(n493), .O(n494));
  nor2   g0422(.a(n413), .b(n85), .O(n495));
  inv1   g0423(.a(n495), .O(n496));
  nor2   g0424(.a(n496), .b(n335), .O(n497));
  nor2   g0425(.a(n339), .b(G77), .O(n498));
  nor2   g0426(.a(n233), .b(n93), .O(n499));
  nor2   g0427(.a(n236), .b(n78), .O(n500));
  nor2   g0428(.a(n85), .b(n83), .O(n501));
  nor2   g0429(.a(n501), .b(n500), .O(n502));
  inv1   g0430(.a(n502), .O(n503));
  nor2   g0431(.a(n503), .b(n499), .O(n504));
  nor2   g0432(.a(n504), .b(n231), .O(n505));
  nor2   g0433(.a(n505), .b(n498), .O(n506));
  inv1   g0434(.a(n506), .O(n507));
  nor2   g0435(.a(n507), .b(n497), .O(n508));
  nor2   g0436(.a(n204), .b(n112), .O(n509));
  nor2   g0437(.a(n207), .b(n94), .O(n510));
  nor2   g0438(.a(n510), .b(n292), .O(n511));
  inv1   g0439(.a(n511), .O(n512));
  nor2   g0440(.a(n512), .b(n509), .O(n513));
  nor2   g0441(.a(n513), .b(n201), .O(n514));
  nor2   g0442(.a(n434), .b(n86), .O(n515));
  nor2   g0443(.a(n515), .b(n432), .O(n516));
  inv1   g0444(.a(n516), .O(n517));
  nor2   g0445(.a(n517), .b(n514), .O(n518));
  nor2   g0446(.a(n518), .b(G169), .O(n519));
  inv1   g0447(.a(n518), .O(n520));
  nor2   g0448(.a(n520), .b(G179), .O(n521));
  nor2   g0449(.a(n521), .b(n519), .O(n522));
  inv1   g0450(.a(n522), .O(n523));
  nor2   g0451(.a(n523), .b(n508), .O(n524));
  nor2   g0452(.a(n518), .b(n260), .O(n525));
  inv1   g0453(.a(n508), .O(n526));
  nor2   g0454(.a(n520), .b(n263), .O(n527));
  nor2   g0455(.a(n527), .b(n526), .O(n528));
  inv1   g0456(.a(n528), .O(n529));
  nor2   g0457(.a(n529), .b(n525), .O(n530));
  nor2   g0458(.a(n530), .b(n524), .O(n531));
  inv1   g0459(.a(n531), .O(n532));
  nor2   g0460(.a(n413), .b(n111), .O(n533));
  inv1   g0461(.a(n533), .O(n534));
  nor2   g0462(.a(n534), .b(n335), .O(n535));
  nor2   g0463(.a(n246), .b(n252), .O(n536));
  nor2   g0464(.a(G68), .b(n83), .O(n537));
  inv1   g0465(.a(n537), .O(n538));
  nor2   g0466(.a(n538), .b(n536), .O(n539));
  nor2   g0467(.a(n233), .b(n106), .O(n540));
  nor2   g0468(.a(n236), .b(n85), .O(n541));
  nor2   g0469(.a(n541), .b(n540), .O(n542));
  nor2   g0470(.a(n542), .b(n231), .O(n543));
  nor2   g0471(.a(n543), .b(n539), .O(n544));
  inv1   g0472(.a(n544), .O(n545));
  nor2   g0473(.a(n545), .b(n535), .O(n546));
  nor2   g0474(.a(n204), .b(n94), .O(n547));
  nor2   g0475(.a(n207), .b(n107), .O(n548));
  nor2   g0476(.a(n96), .b(n197), .O(n549));
  nor2   g0477(.a(n549), .b(n548), .O(n550));
  inv1   g0478(.a(n550), .O(n551));
  nor2   g0479(.a(n551), .b(n547), .O(n552));
  nor2   g0480(.a(n552), .b(n201), .O(n553));
  nor2   g0481(.a(n434), .b(n112), .O(n554));
  nor2   g0482(.a(n554), .b(n432), .O(n555));
  inv1   g0483(.a(n555), .O(n556));
  nor2   g0484(.a(n556), .b(n553), .O(n557));
  nor2   g0485(.a(n557), .b(G169), .O(n558));
  inv1   g0486(.a(n557), .O(n559));
  nor2   g0487(.a(n559), .b(G179), .O(n560));
  nor2   g0488(.a(n560), .b(n558), .O(n561));
  inv1   g0489(.a(n561), .O(n562));
  nor2   g0490(.a(n562), .b(n546), .O(n563));
  nor2   g0491(.a(n557), .b(n260), .O(n564));
  inv1   g0492(.a(n546), .O(n565));
  nor2   g0493(.a(n559), .b(n263), .O(n566));
  nor2   g0494(.a(n566), .b(n565), .O(n567));
  inv1   g0495(.a(n567), .O(n568));
  nor2   g0496(.a(n568), .b(n564), .O(n569));
  nor2   g0497(.a(n569), .b(n563), .O(n570));
  inv1   g0498(.a(n570), .O(n571));
  nor2   g0499(.a(n571), .b(n532), .O(n572));
  inv1   g0500(.a(n572), .O(n573));
  nor2   g0501(.a(n573), .b(n494), .O(n574));
  inv1   g0502(.a(n574), .O(n575));
  nor2   g0503(.a(n575), .b(n403), .O(G372));
  inv1   g0504(.a(n351), .O(n577));
  nor2   g0505(.a(n397), .b(n577), .O(n578));
  nor2   g0506(.a(n578), .b(n391), .O(n579));
  nor2   g0507(.a(n579), .b(n316), .O(n580));
  inv1   g0508(.a(n306), .O(n581));
  nor2   g0509(.a(n581), .b(n267), .O(n582));
  nor2   g0510(.a(n582), .b(n259), .O(n583));
  inv1   g0511(.a(n583), .O(n584));
  nor2   g0512(.a(n584), .b(n580), .O(n585));
  nor2   g0513(.a(n585), .b(n575), .O(n586));
  inv1   g0514(.a(n524), .O(n587));
  nor2   g0515(.a(n569), .b(n587), .O(n588));
  nor2   g0516(.a(n588), .b(n563), .O(n589));
  nor2   g0517(.a(n589), .b(n494), .O(n590));
  inv1   g0518(.a(n484), .O(n591));
  nor2   g0519(.a(n591), .b(n450), .O(n592));
  nor2   g0520(.a(n592), .b(n444), .O(n593));
  inv1   g0521(.a(n593), .O(n594));
  nor2   g0522(.a(n594), .b(n590), .O(n595));
  inv1   g0523(.a(n595), .O(n596));
  nor2   g0524(.a(n596), .b(n586), .O(n597));
  inv1   g0525(.a(n597), .O(G369));
  inv1   g0526(.a(n391), .O(n599));
  inv1   g0527(.a(G343), .O(n600));
  inv1   g0528(.a(G213), .O(n601));
  nor2   g0529(.a(n601), .b(G20), .O(n602));
  inv1   g0530(.a(n602), .O(n603));
  nor2   g0531(.a(n603), .b(n247), .O(n604));
  inv1   g0532(.a(n604), .O(n605));
  nor2   g0533(.a(n605), .b(n600), .O(n606));
  nor2   g0534(.a(n606), .b(n599), .O(n607));
  nor2   g0535(.a(n606), .b(n577), .O(n608));
  inv1   g0536(.a(n608), .O(n609));
  inv1   g0537(.a(n606), .O(n610));
  nor2   g0538(.a(n610), .b(n373), .O(n611));
  nor2   g0539(.a(n611), .b(n399), .O(n612));
  inv1   g0540(.a(n611), .O(n613));
  nor2   g0541(.a(n613), .b(n599), .O(n614));
  nor2   g0542(.a(n614), .b(n612), .O(n615));
  nor2   g0543(.a(n615), .b(n609), .O(n616));
  nor2   g0544(.a(n616), .b(n607), .O(n617));
  inv1   g0545(.a(n617), .O(n618));
  inv1   g0546(.a(G330), .O(n619));
  nor2   g0547(.a(n610), .b(n350), .O(n620));
  nor2   g0548(.a(n620), .b(n359), .O(n621));
  nor2   g0549(.a(n610), .b(n577), .O(n622));
  nor2   g0550(.a(n622), .b(n621), .O(n623));
  nor2   g0551(.a(n623), .b(n619), .O(n624));
  inv1   g0552(.a(n624), .O(n625));
  nor2   g0553(.a(n625), .b(n615), .O(n626));
  nor2   g0554(.a(n626), .b(n618), .O(n627));
  inv1   g0555(.a(n627), .O(G399));
  nor2   g0556(.a(n606), .b(n585), .O(n629));
  inv1   g0557(.a(n333), .O(n630));
  nor2   g0558(.a(n387), .b(n226), .O(n631));
  inv1   g0559(.a(n631), .O(n632));
  nor2   g0560(.a(n632), .b(n287), .O(n633));
  inv1   g0561(.a(n633), .O(n634));
  nor2   g0562(.a(n634), .b(n630), .O(n635));
  nor2   g0563(.a(n329), .b(G179), .O(n636));
  inv1   g0564(.a(n636), .O(n637));
  nor2   g0565(.a(n385), .b(n225), .O(n638));
  inv1   g0566(.a(n638), .O(n639));
  nor2   g0567(.a(n639), .b(n286), .O(n640));
  inv1   g0568(.a(n640), .O(n641));
  nor2   g0569(.a(n641), .b(n637), .O(n642));
  nor2   g0570(.a(n642), .b(n635), .O(n643));
  nor2   g0571(.a(n643), .b(n610), .O(n644));
  nor2   g0572(.a(n606), .b(n403), .O(n645));
  nor2   g0573(.a(n645), .b(n644), .O(n646));
  nor2   g0574(.a(n646), .b(n619), .O(n647));
  nor2   g0575(.a(n647), .b(n629), .O(n648));
  nor2   g0576(.a(n648), .b(G1), .O(n649));
  nor2   g0577(.a(n134), .b(G41), .O(n650));
  inv1   g0578(.a(n240), .O(n651));
  nor2   g0579(.a(n651), .b(G116), .O(n652));
  inv1   g0580(.a(n652), .O(n653));
  nor2   g0581(.a(n653), .b(n82), .O(n654));
  inv1   g0582(.a(n654), .O(n655));
  nor2   g0583(.a(n655), .b(n650), .O(n656));
  inv1   g0584(.a(n650), .O(n657));
  nor2   g0585(.a(n657), .b(n129), .O(n658));
  nor2   g0586(.a(n658), .b(n656), .O(n659));
  inv1   g0587(.a(n659), .O(n660));
  nor2   g0588(.a(n660), .b(n649), .O(n661));
  inv1   g0589(.a(n661), .O(G364));
  inv1   g0590(.a(n623), .O(n663));
  nor2   g0591(.a(G20), .b(G13), .O(n664));
  inv1   g0592(.a(n664), .O(n665));
  nor2   g0593(.a(n665), .b(G33), .O(n666));
  inv1   g0594(.a(n666), .O(n667));
  nor2   g0595(.a(n667), .b(n663), .O(n668));
  nor2   g0596(.a(G169), .b(n83), .O(n669));
  nor2   g0597(.a(n669), .b(n124), .O(n670));
  nor2   g0598(.a(n670), .b(n666), .O(n671));
  inv1   g0599(.a(n671), .O(n672));
  nor2   g0600(.a(n192), .b(n216), .O(n673));
  nor2   g0601(.a(n134), .b(n197), .O(n674));
  inv1   g0602(.a(n674), .O(n675));
  nor2   g0603(.a(n129), .b(G45), .O(n676));
  nor2   g0604(.a(n676), .b(n675), .O(n677));
  inv1   g0605(.a(n677), .O(n678));
  nor2   g0606(.a(n678), .b(n673), .O(n679));
  nor2   g0607(.a(n133), .b(G116), .O(n680));
  nor2   g0608(.a(n134), .b(G33), .O(n681));
  inv1   g0609(.a(n681), .O(n682));
  nor2   g0610(.a(n682), .b(n80), .O(n683));
  nor2   g0611(.a(n683), .b(n680), .O(n684));
  inv1   g0612(.a(n684), .O(n685));
  nor2   g0613(.a(n685), .b(n679), .O(n686));
  nor2   g0614(.a(n686), .b(n672), .O(n687));
  nor2   g0615(.a(G20), .b(n122), .O(n688));
  inv1   g0616(.a(n688), .O(n689));
  nor2   g0617(.a(n689), .b(n216), .O(n690));
  nor2   g0618(.a(n690), .b(n82), .O(n691));
  inv1   g0619(.a(n691), .O(n692));
  nor2   g0620(.a(n692), .b(n650), .O(n693));
  inv1   g0621(.a(n693), .O(n694));
  inv1   g0622(.a(n670), .O(n695));
  nor2   g0623(.a(n331), .b(n83), .O(n696));
  nor2   g0624(.a(n260), .b(n83), .O(n697));
  inv1   g0625(.a(n697), .O(n698));
  nor2   g0626(.a(n698), .b(n696), .O(n699));
  inv1   g0627(.a(n699), .O(n700));
  nor2   g0628(.a(n700), .b(G190), .O(n701));
  inv1   g0629(.a(n701), .O(n702));
  nor2   g0630(.a(n702), .b(n103), .O(n703));
  nor2   g0631(.a(G190), .b(n83), .O(n704));
  nor2   g0632(.a(n697), .b(n696), .O(n705));
  inv1   g0633(.a(n705), .O(n706));
  nor2   g0634(.a(n706), .b(n704), .O(n707));
  inv1   g0635(.a(n707), .O(n708));
  nor2   g0636(.a(n708), .b(n96), .O(n709));
  inv1   g0637(.a(n704), .O(n710));
  nor2   g0638(.a(n706), .b(n710), .O(n711));
  inv1   g0639(.a(n711), .O(n712));
  nor2   g0640(.a(n712), .b(n453), .O(n713));
  nor2   g0641(.a(n713), .b(n709), .O(n714));
  inv1   g0642(.a(n714), .O(n715));
  nor2   g0643(.a(n715), .b(n703), .O(n716));
  inv1   g0644(.a(n716), .O(n717));
  inv1   g0645(.a(n696), .O(n718));
  nor2   g0646(.a(n718), .b(n260), .O(n719));
  inv1   g0647(.a(n719), .O(n720));
  nor2   g0648(.a(n720), .b(n263), .O(n721));
  inv1   g0649(.a(n721), .O(n722));
  nor2   g0650(.a(n722), .b(n106), .O(n723));
  nor2   g0651(.a(n723), .b(G33), .O(n724));
  inv1   g0652(.a(n724), .O(n725));
  nor2   g0653(.a(n720), .b(G190), .O(n726));
  inv1   g0654(.a(n726), .O(n727));
  nor2   g0655(.a(n727), .b(n111), .O(n728));
  nor2   g0656(.a(n718), .b(G200), .O(n729));
  inv1   g0657(.a(n729), .O(n730));
  nor2   g0658(.a(n730), .b(n263), .O(n731));
  inv1   g0659(.a(n731), .O(n732));
  nor2   g0660(.a(n732), .b(n93), .O(n733));
  nor2   g0661(.a(n733), .b(n728), .O(n734));
  inv1   g0662(.a(n734), .O(n735));
  nor2   g0663(.a(n730), .b(G190), .O(n736));
  inv1   g0664(.a(n736), .O(n737));
  nor2   g0665(.a(n737), .b(n85), .O(n738));
  nor2   g0666(.a(n700), .b(n263), .O(n739));
  inv1   g0667(.a(n739), .O(n740));
  nor2   g0668(.a(n740), .b(n78), .O(n741));
  nor2   g0669(.a(n741), .b(n738), .O(n742));
  inv1   g0670(.a(n742), .O(n743));
  nor2   g0671(.a(n743), .b(n735), .O(n744));
  inv1   g0672(.a(n744), .O(n745));
  nor2   g0673(.a(n745), .b(n725), .O(n746));
  inv1   g0674(.a(n746), .O(n747));
  nor2   g0675(.a(n747), .b(n717), .O(n748));
  nor2   g0676(.a(n702), .b(n272), .O(n749));
  inv1   g0677(.a(G329), .O(n750));
  nor2   g0678(.a(n712), .b(n750), .O(n751));
  nor2   g0679(.a(n708), .b(n375), .O(n752));
  nor2   g0680(.a(n752), .b(n751), .O(n753));
  inv1   g0681(.a(n753), .O(n754));
  nor2   g0682(.a(n754), .b(n749), .O(n755));
  inv1   g0683(.a(n755), .O(n756));
  inv1   g0684(.a(G326), .O(n757));
  nor2   g0685(.a(n722), .b(n757), .O(n758));
  nor2   g0686(.a(n758), .b(n197), .O(n759));
  inv1   g0687(.a(n759), .O(n760));
  inv1   g0688(.a(G317), .O(n761));
  nor2   g0689(.a(n727), .b(n761), .O(n762));
  inv1   g0690(.a(G322), .O(n763));
  nor2   g0691(.a(n732), .b(n763), .O(n764));
  nor2   g0692(.a(n764), .b(n762), .O(n765));
  inv1   g0693(.a(n765), .O(n766));
  inv1   g0694(.a(G311), .O(n767));
  nor2   g0695(.a(n737), .b(n767), .O(n768));
  nor2   g0696(.a(n740), .b(n320), .O(n769));
  nor2   g0697(.a(n769), .b(n768), .O(n770));
  inv1   g0698(.a(n770), .O(n771));
  nor2   g0699(.a(n771), .b(n766), .O(n772));
  inv1   g0700(.a(n772), .O(n773));
  nor2   g0701(.a(n773), .b(n760), .O(n774));
  inv1   g0702(.a(n774), .O(n775));
  nor2   g0703(.a(n775), .b(n756), .O(n776));
  nor2   g0704(.a(n776), .b(n748), .O(n777));
  nor2   g0705(.a(n777), .b(n695), .O(n778));
  nor2   g0706(.a(n778), .b(n694), .O(n779));
  inv1   g0707(.a(n779), .O(n780));
  nor2   g0708(.a(n780), .b(n687), .O(n781));
  inv1   g0709(.a(n781), .O(n782));
  nor2   g0710(.a(n782), .b(n668), .O(n783));
  nor2   g0711(.a(n663), .b(G330), .O(n784));
  nor2   g0712(.a(n693), .b(n624), .O(n785));
  inv1   g0713(.a(n785), .O(n786));
  nor2   g0714(.a(n786), .b(n784), .O(n787));
  nor2   g0715(.a(n787), .b(n783), .O(n788));
  inv1   g0716(.a(n788), .O(G396));
  nor2   g0717(.a(G33), .b(G13), .O(n790));
  inv1   g0718(.a(n790), .O(n791));
  nor2   g0719(.a(n610), .b(n508), .O(n792));
  nor2   g0720(.a(n792), .b(n532), .O(n793));
  inv1   g0721(.a(n792), .O(n794));
  nor2   g0722(.a(n794), .b(n587), .O(n795));
  nor2   g0723(.a(n795), .b(n793), .O(n796));
  inv1   g0724(.a(n796), .O(n797));
  nor2   g0725(.a(n797), .b(n791), .O(n798));
  nor2   g0726(.a(n702), .b(n111), .O(n799));
  nor2   g0727(.a(n708), .b(n93), .O(n800));
  inv1   g0728(.a(G132), .O(n801));
  nor2   g0729(.a(n712), .b(n801), .O(n802));
  nor2   g0730(.a(n802), .b(n800), .O(n803));
  inv1   g0731(.a(n803), .O(n804));
  nor2   g0732(.a(n804), .b(n799), .O(n805));
  inv1   g0733(.a(n805), .O(n806));
  inv1   g0734(.a(G137), .O(n807));
  nor2   g0735(.a(n722), .b(n807), .O(n808));
  nor2   g0736(.a(n808), .b(G33), .O(n809));
  inv1   g0737(.a(n809), .O(n810));
  nor2   g0738(.a(n727), .b(n404), .O(n811));
  inv1   g0739(.a(G143), .O(n812));
  nor2   g0740(.a(n732), .b(n812), .O(n813));
  nor2   g0741(.a(n813), .b(n811), .O(n814));
  inv1   g0742(.a(n814), .O(n815));
  nor2   g0743(.a(n737), .b(n453), .O(n816));
  nor2   g0744(.a(n740), .b(n106), .O(n817));
  nor2   g0745(.a(n817), .b(n816), .O(n818));
  inv1   g0746(.a(n818), .O(n819));
  nor2   g0747(.a(n819), .b(n815), .O(n820));
  inv1   g0748(.a(n820), .O(n821));
  nor2   g0749(.a(n821), .b(n810), .O(n822));
  inv1   g0750(.a(n822), .O(n823));
  nor2   g0751(.a(n823), .b(n806), .O(n824));
  nor2   g0752(.a(n712), .b(n767), .O(n825));
  nor2   g0753(.a(n702), .b(n78), .O(n826));
  nor2   g0754(.a(n737), .b(n88), .O(n827));
  nor2   g0755(.a(n827), .b(n826), .O(n828));
  inv1   g0756(.a(n828), .O(n829));
  nor2   g0757(.a(n829), .b(n825), .O(n830));
  inv1   g0758(.a(n830), .O(n831));
  nor2   g0759(.a(n709), .b(n197), .O(n832));
  inv1   g0760(.a(n832), .O(n833));
  nor2   g0761(.a(n740), .b(n103), .O(n834));
  nor2   g0762(.a(n732), .b(n375), .O(n835));
  nor2   g0763(.a(n835), .b(n834), .O(n836));
  inv1   g0764(.a(n836), .O(n837));
  nor2   g0765(.a(n722), .b(n320), .O(n838));
  nor2   g0766(.a(n727), .b(n272), .O(n839));
  nor2   g0767(.a(n839), .b(n838), .O(n840));
  inv1   g0768(.a(n840), .O(n841));
  nor2   g0769(.a(n841), .b(n837), .O(n842));
  inv1   g0770(.a(n842), .O(n843));
  nor2   g0771(.a(n843), .b(n833), .O(n844));
  inv1   g0772(.a(n844), .O(n845));
  nor2   g0773(.a(n845), .b(n831), .O(n846));
  nor2   g0774(.a(n846), .b(n824), .O(n847));
  nor2   g0775(.a(n847), .b(n695), .O(n848));
  nor2   g0776(.a(n790), .b(n670), .O(n849));
  inv1   g0777(.a(n849), .O(n850));
  nor2   g0778(.a(n850), .b(G77), .O(n851));
  nor2   g0779(.a(n851), .b(n694), .O(n852));
  inv1   g0780(.a(n852), .O(n853));
  nor2   g0781(.a(n853), .b(n848), .O(n854));
  inv1   g0782(.a(n854), .O(n855));
  nor2   g0783(.a(n855), .b(n798), .O(n856));
  inv1   g0784(.a(n647), .O(n857));
  inv1   g0785(.a(n629), .O(n858));
  nor2   g0786(.a(n796), .b(n858), .O(n859));
  nor2   g0787(.a(n797), .b(n629), .O(n860));
  nor2   g0788(.a(n860), .b(n859), .O(n861));
  inv1   g0789(.a(n861), .O(n862));
  nor2   g0790(.a(n862), .b(n857), .O(n863));
  nor2   g0791(.a(n861), .b(n647), .O(n864));
  nor2   g0792(.a(n864), .b(n693), .O(n865));
  inv1   g0793(.a(n865), .O(n866));
  nor2   g0794(.a(n866), .b(n863), .O(n867));
  nor2   g0795(.a(n867), .b(n856), .O(n868));
  inv1   g0796(.a(n868), .O(G384));
  nor2   g0797(.a(n604), .b(n591), .O(n870));
  inv1   g0798(.a(n563), .O(n871));
  nor2   g0799(.a(n606), .b(n871), .O(n872));
  nor2   g0800(.a(n606), .b(n587), .O(n873));
  nor2   g0801(.a(n873), .b(n859), .O(n874));
  nor2   g0802(.a(n610), .b(n546), .O(n875));
  nor2   g0803(.a(n875), .b(n571), .O(n876));
  inv1   g0804(.a(n875), .O(n877));
  nor2   g0805(.a(n877), .b(n871), .O(n878));
  nor2   g0806(.a(n878), .b(n876), .O(n879));
  nor2   g0807(.a(n879), .b(n874), .O(n880));
  nor2   g0808(.a(n880), .b(n872), .O(n881));
  nor2   g0809(.a(n605), .b(n467), .O(n882));
  nor2   g0810(.a(n882), .b(n492), .O(n883));
  inv1   g0811(.a(n882), .O(n884));
  nor2   g0812(.a(n884), .b(n591), .O(n885));
  nor2   g0813(.a(n885), .b(n883), .O(n886));
  nor2   g0814(.a(n886), .b(n881), .O(n887));
  nor2   g0815(.a(n887), .b(n870), .O(n888));
  nor2   g0816(.a(n879), .b(n796), .O(n889));
  inv1   g0817(.a(n889), .O(n890));
  nor2   g0818(.a(n890), .b(n886), .O(n891));
  nor2   g0819(.a(n891), .b(n646), .O(n892));
  nor2   g0820(.a(n892), .b(n575), .O(n893));
  inv1   g0821(.a(n891), .O(n894));
  nor2   g0822(.a(n894), .b(n646), .O(n895));
  nor2   g0823(.a(n895), .b(n574), .O(n896));
  nor2   g0824(.a(n896), .b(n619), .O(n897));
  inv1   g0825(.a(n897), .O(n898));
  nor2   g0826(.a(n898), .b(n893), .O(n899));
  nor2   g0827(.a(n899), .b(n888), .O(n900));
  inv1   g0828(.a(n888), .O(n901));
  inv1   g0829(.a(n899), .O(n902));
  nor2   g0830(.a(n902), .b(n901), .O(n903));
  nor2   g0831(.a(n903), .b(n900), .O(n904));
  inv1   g0832(.a(n904), .O(n905));
  nor2   g0833(.a(n858), .b(n575), .O(n906));
  nor2   g0834(.a(n906), .b(n596), .O(n907));
  inv1   g0835(.a(n907), .O(n908));
  nor2   g0836(.a(n908), .b(n905), .O(n909));
  nor2   g0837(.a(n907), .b(n904), .O(n910));
  nor2   g0838(.a(n131), .b(n125), .O(n911));
  inv1   g0839(.a(n911), .O(n912));
  nor2   g0840(.a(n912), .b(n910), .O(n913));
  inv1   g0841(.a(n913), .O(n914));
  nor2   g0842(.a(n914), .b(n909), .O(n915));
  nor2   g0843(.a(n185), .b(n106), .O(n916));
  nor2   g0844(.a(G68), .b(G50), .O(n917));
  nor2   g0845(.a(n917), .b(n132), .O(n918));
  inv1   g0846(.a(n918), .O(n919));
  nor2   g0847(.a(n919), .b(n916), .O(n920));
  nor2   g0848(.a(n126), .b(n88), .O(n921));
  inv1   g0849(.a(n921), .O(n922));
  nor2   g0850(.a(n922), .b(n172), .O(n923));
  nor2   g0851(.a(n923), .b(n920), .O(n924));
  inv1   g0852(.a(n924), .O(n925));
  nor2   g0853(.a(n925), .b(n915), .O(n926));
  inv1   g0854(.a(n926), .O(G367));
  inv1   g0855(.a(n648), .O(n928));
  inv1   g0856(.a(n615), .O(n929));
  nor2   g0857(.a(n929), .b(n608), .O(n930));
  nor2   g0858(.a(n930), .b(n616), .O(n931));
  inv1   g0859(.a(n931), .O(n932));
  nor2   g0860(.a(n932), .b(n625), .O(n933));
  nor2   g0861(.a(n931), .b(n624), .O(n934));
  nor2   g0862(.a(n934), .b(n933), .O(n935));
  inv1   g0863(.a(n935), .O(n936));
  nor2   g0864(.a(n936), .b(n928), .O(n937));
  inv1   g0865(.a(n937), .O(n938));
  nor2   g0866(.a(n610), .b(n303), .O(n939));
  nor2   g0867(.a(n939), .b(n314), .O(n940));
  inv1   g0868(.a(n939), .O(n941));
  nor2   g0869(.a(n941), .b(n581), .O(n942));
  nor2   g0870(.a(n942), .b(n940), .O(n943));
  inv1   g0871(.a(n943), .O(n944));
  inv1   g0872(.a(n626), .O(n945));
  nor2   g0873(.a(n945), .b(n617), .O(n946));
  nor2   g0874(.a(n946), .b(n627), .O(n947));
  inv1   g0875(.a(n947), .O(n948));
  nor2   g0876(.a(n948), .b(n944), .O(n949));
  nor2   g0877(.a(n947), .b(n943), .O(n950));
  nor2   g0878(.a(n950), .b(n949), .O(n951));
  nor2   g0879(.a(n951), .b(n938), .O(n952));
  nor2   g0880(.a(n952), .b(n928), .O(n953));
  nor2   g0881(.a(n606), .b(n581), .O(n954));
  nor2   g0882(.a(n943), .b(n617), .O(n955));
  nor2   g0883(.a(n955), .b(n954), .O(n956));
  inv1   g0884(.a(n956), .O(n957));
  nor2   g0885(.a(n943), .b(n945), .O(n958));
  nor2   g0886(.a(n958), .b(n957), .O(n959));
  inv1   g0887(.a(n958), .O(n960));
  nor2   g0888(.a(n960), .b(n956), .O(n961));
  nor2   g0889(.a(n961), .b(n959), .O(n962));
  inv1   g0890(.a(n962), .O(n963));
  nor2   g0891(.a(n610), .b(n256), .O(n964));
  nor2   g0892(.a(n964), .b(n269), .O(n965));
  inv1   g0893(.a(n259), .O(n966));
  inv1   g0894(.a(n964), .O(n967));
  nor2   g0895(.a(n967), .b(n966), .O(n968));
  nor2   g0896(.a(n968), .b(n965), .O(n969));
  inv1   g0897(.a(n969), .O(n970));
  nor2   g0898(.a(n970), .b(n963), .O(n971));
  nor2   g0899(.a(n969), .b(n962), .O(n972));
  nor2   g0900(.a(n972), .b(n971), .O(n973));
  nor2   g0901(.a(n973), .b(n657), .O(n974));
  inv1   g0902(.a(n974), .O(n975));
  nor2   g0903(.a(n975), .b(n953), .O(n976));
  nor2   g0904(.a(n973), .b(n691), .O(n977));
  nor2   g0905(.a(n970), .b(n667), .O(n978));
  nor2   g0906(.a(n702), .b(n85), .O(n979));
  nor2   g0907(.a(n708), .b(n111), .O(n980));
  nor2   g0908(.a(n712), .b(n807), .O(n981));
  nor2   g0909(.a(n981), .b(n980), .O(n982));
  inv1   g0910(.a(n982), .O(n983));
  nor2   g0911(.a(n983), .b(n979), .O(n984));
  inv1   g0912(.a(n984), .O(n985));
  nor2   g0913(.a(n722), .b(n812), .O(n986));
  nor2   g0914(.a(n986), .b(G33), .O(n987));
  inv1   g0915(.a(n987), .O(n988));
  nor2   g0916(.a(n727), .b(n453), .O(n989));
  nor2   g0917(.a(n732), .b(n404), .O(n990));
  nor2   g0918(.a(n990), .b(n989), .O(n991));
  inv1   g0919(.a(n991), .O(n992));
  nor2   g0920(.a(n737), .b(n106), .O(n993));
  nor2   g0921(.a(n740), .b(n93), .O(n994));
  nor2   g0922(.a(n994), .b(n993), .O(n995));
  inv1   g0923(.a(n995), .O(n996));
  nor2   g0924(.a(n996), .b(n992), .O(n997));
  inv1   g0925(.a(n997), .O(n998));
  nor2   g0926(.a(n998), .b(n988), .O(n999));
  inv1   g0927(.a(n999), .O(n1000));
  nor2   g0928(.a(n1000), .b(n985), .O(n1001));
  nor2   g0929(.a(n702), .b(n96), .O(n1002));
  nor2   g0930(.a(n708), .b(n103), .O(n1003));
  nor2   g0931(.a(n712), .b(n761), .O(n1004));
  nor2   g0932(.a(n1004), .b(n1003), .O(n1005));
  inv1   g0933(.a(n1005), .O(n1006));
  nor2   g0934(.a(n1006), .b(n1002), .O(n1007));
  inv1   g0935(.a(n1007), .O(n1008));
  nor2   g0936(.a(n722), .b(n767), .O(n1009));
  nor2   g0937(.a(n1009), .b(n197), .O(n1010));
  inv1   g0938(.a(n1010), .O(n1011));
  nor2   g0939(.a(n727), .b(n375), .O(n1012));
  nor2   g0940(.a(n732), .b(n320), .O(n1013));
  nor2   g0941(.a(n1013), .b(n1012), .O(n1014));
  inv1   g0942(.a(n1014), .O(n1015));
  nor2   g0943(.a(n737), .b(n272), .O(n1016));
  nor2   g0944(.a(n740), .b(n88), .O(n1017));
  nor2   g0945(.a(n1017), .b(n1016), .O(n1018));
  inv1   g0946(.a(n1018), .O(n1019));
  nor2   g0947(.a(n1019), .b(n1015), .O(n1020));
  inv1   g0948(.a(n1020), .O(n1021));
  nor2   g0949(.a(n1021), .b(n1011), .O(n1022));
  inv1   g0950(.a(n1022), .O(n1023));
  nor2   g0951(.a(n1023), .b(n1008), .O(n1024));
  nor2   g0952(.a(n1024), .b(n1001), .O(n1025));
  nor2   g0953(.a(n1025), .b(n695), .O(n1026));
  nor2   g0954(.a(n675), .b(n153), .O(n1027));
  nor2   g0955(.a(n133), .b(G87), .O(n1028));
  nor2   g0956(.a(n1028), .b(n681), .O(n1029));
  inv1   g0957(.a(n1029), .O(n1030));
  nor2   g0958(.a(n1030), .b(n1027), .O(n1031));
  nor2   g0959(.a(n1031), .b(n672), .O(n1032));
  nor2   g0960(.a(n1032), .b(n694), .O(n1033));
  inv1   g0961(.a(n1033), .O(n1034));
  nor2   g0962(.a(n1034), .b(n1026), .O(n1035));
  inv1   g0963(.a(n1035), .O(n1036));
  nor2   g0964(.a(n1036), .b(n978), .O(n1037));
  nor2   g0965(.a(n1037), .b(n977), .O(n1038));
  inv1   g0966(.a(n1038), .O(n1039));
  nor2   g0967(.a(n1039), .b(n976), .O(n1040));
  inv1   g0968(.a(n1040), .O(G387));
  nor2   g0969(.a(n935), .b(n648), .O(n1042));
  nor2   g0970(.a(n937), .b(n657), .O(n1043));
  inv1   g0971(.a(n1043), .O(n1044));
  nor2   g0972(.a(n1044), .b(n1042), .O(n1045));
  nor2   g0973(.a(n936), .b(n691), .O(n1046));
  nor2   g0974(.a(n667), .b(n929), .O(n1047));
  nor2   g0975(.a(n164), .b(n216), .O(n1048));
  nor2   g0976(.a(n85), .b(n111), .O(n1049));
  nor2   g0977(.a(G50), .b(G45), .O(n1050));
  inv1   g0978(.a(n1050), .O(n1051));
  nor2   g0979(.a(n1051), .b(n93), .O(n1052));
  inv1   g0980(.a(n1052), .O(n1053));
  nor2   g0981(.a(n1053), .b(n1049), .O(n1054));
  inv1   g0982(.a(n1054), .O(n1055));
  nor2   g0983(.a(n1055), .b(n653), .O(n1056));
  nor2   g0984(.a(n1056), .b(n675), .O(n1057));
  inv1   g0985(.a(n1057), .O(n1058));
  nor2   g0986(.a(n1058), .b(n1048), .O(n1059));
  nor2   g0987(.a(n133), .b(G107), .O(n1060));
  nor2   g0988(.a(n682), .b(n652), .O(n1061));
  nor2   g0989(.a(n1061), .b(n1060), .O(n1062));
  inv1   g0990(.a(n1062), .O(n1063));
  nor2   g0991(.a(n1063), .b(n1059), .O(n1064));
  nor2   g0992(.a(n1064), .b(n672), .O(n1065));
  nor2   g0993(.a(n708), .b(n78), .O(n1066));
  nor2   g0994(.a(n712), .b(n404), .O(n1067));
  nor2   g0995(.a(n737), .b(n111), .O(n1068));
  nor2   g0996(.a(n1068), .b(n1067), .O(n1069));
  inv1   g0997(.a(n1069), .O(n1070));
  nor2   g0998(.a(n1070), .b(n1066), .O(n1071));
  inv1   g0999(.a(n1071), .O(n1072));
  nor2   g1000(.a(n1002), .b(G33), .O(n1073));
  inv1   g1001(.a(n1073), .O(n1074));
  nor2   g1002(.a(n740), .b(n85), .O(n1075));
  nor2   g1003(.a(n732), .b(n106), .O(n1076));
  nor2   g1004(.a(n1076), .b(n1075), .O(n1077));
  inv1   g1005(.a(n1077), .O(n1078));
  nor2   g1006(.a(n722), .b(n453), .O(n1079));
  nor2   g1007(.a(n727), .b(n93), .O(n1080));
  nor2   g1008(.a(n1080), .b(n1079), .O(n1081));
  inv1   g1009(.a(n1081), .O(n1082));
  nor2   g1010(.a(n1082), .b(n1078), .O(n1083));
  inv1   g1011(.a(n1083), .O(n1084));
  nor2   g1012(.a(n1084), .b(n1074), .O(n1085));
  inv1   g1013(.a(n1085), .O(n1086));
  nor2   g1014(.a(n1086), .b(n1072), .O(n1087));
  nor2   g1015(.a(n702), .b(n88), .O(n1088));
  nor2   g1016(.a(n708), .b(n272), .O(n1089));
  nor2   g1017(.a(n712), .b(n757), .O(n1090));
  nor2   g1018(.a(n1090), .b(n1089), .O(n1091));
  inv1   g1019(.a(n1091), .O(n1092));
  nor2   g1020(.a(n1092), .b(n1088), .O(n1093));
  inv1   g1021(.a(n1093), .O(n1094));
  nor2   g1022(.a(n722), .b(n763), .O(n1095));
  nor2   g1023(.a(n1095), .b(n197), .O(n1096));
  inv1   g1024(.a(n1096), .O(n1097));
  nor2   g1025(.a(n727), .b(n767), .O(n1098));
  nor2   g1026(.a(n732), .b(n761), .O(n1099));
  nor2   g1027(.a(n1099), .b(n1098), .O(n1100));
  inv1   g1028(.a(n1100), .O(n1101));
  nor2   g1029(.a(n737), .b(n320), .O(n1102));
  nor2   g1030(.a(n740), .b(n375), .O(n1103));
  nor2   g1031(.a(n1103), .b(n1102), .O(n1104));
  inv1   g1032(.a(n1104), .O(n1105));
  nor2   g1033(.a(n1105), .b(n1101), .O(n1106));
  inv1   g1034(.a(n1106), .O(n1107));
  nor2   g1035(.a(n1107), .b(n1097), .O(n1108));
  inv1   g1036(.a(n1108), .O(n1109));
  nor2   g1037(.a(n1109), .b(n1094), .O(n1110));
  nor2   g1038(.a(n1110), .b(n1087), .O(n1111));
  nor2   g1039(.a(n1111), .b(n695), .O(n1112));
  nor2   g1040(.a(n1112), .b(n694), .O(n1113));
  inv1   g1041(.a(n1113), .O(n1114));
  nor2   g1042(.a(n1114), .b(n1065), .O(n1115));
  inv1   g1043(.a(n1115), .O(n1116));
  nor2   g1044(.a(n1116), .b(n1047), .O(n1117));
  nor2   g1045(.a(n1117), .b(n1046), .O(n1118));
  inv1   g1046(.a(n1118), .O(n1119));
  nor2   g1047(.a(n1119), .b(n1045), .O(n1120));
  inv1   g1048(.a(n1120), .O(G393));
  inv1   g1049(.a(n951), .O(n1122));
  nor2   g1050(.a(n1122), .b(n937), .O(n1123));
  nor2   g1051(.a(n952), .b(n657), .O(n1124));
  inv1   g1052(.a(n1124), .O(n1125));
  nor2   g1053(.a(n1125), .b(n1123), .O(n1126));
  nor2   g1054(.a(n951), .b(n691), .O(n1127));
  nor2   g1055(.a(n944), .b(n667), .O(n1128));
  nor2   g1056(.a(n708), .b(n85), .O(n1129));
  nor2   g1057(.a(n712), .b(n812), .O(n1130));
  nor2   g1058(.a(n737), .b(n93), .O(n1131));
  nor2   g1059(.a(n1131), .b(n1130), .O(n1132));
  inv1   g1060(.a(n1132), .O(n1133));
  nor2   g1061(.a(n1133), .b(n1129), .O(n1134));
  inv1   g1062(.a(n1134), .O(n1135));
  nor2   g1063(.a(n826), .b(G33), .O(n1136));
  inv1   g1064(.a(n1136), .O(n1137));
  nor2   g1065(.a(n740), .b(n111), .O(n1138));
  nor2   g1066(.a(n732), .b(n453), .O(n1139));
  nor2   g1067(.a(n1139), .b(n1138), .O(n1140));
  inv1   g1068(.a(n1140), .O(n1141));
  nor2   g1069(.a(n722), .b(n404), .O(n1142));
  nor2   g1070(.a(n727), .b(n106), .O(n1143));
  nor2   g1071(.a(n1143), .b(n1142), .O(n1144));
  inv1   g1072(.a(n1144), .O(n1145));
  nor2   g1073(.a(n1145), .b(n1141), .O(n1146));
  inv1   g1074(.a(n1146), .O(n1147));
  nor2   g1075(.a(n1147), .b(n1137), .O(n1148));
  inv1   g1076(.a(n1148), .O(n1149));
  nor2   g1077(.a(n1149), .b(n1135), .O(n1150));
  nor2   g1078(.a(n708), .b(n88), .O(n1151));
  nor2   g1079(.a(n712), .b(n763), .O(n1152));
  nor2   g1080(.a(n737), .b(n375), .O(n1153));
  nor2   g1081(.a(n1153), .b(n1152), .O(n1154));
  inv1   g1082(.a(n1154), .O(n1155));
  nor2   g1083(.a(n1155), .b(n1151), .O(n1156));
  inv1   g1084(.a(n1156), .O(n1157));
  nor2   g1085(.a(n703), .b(n197), .O(n1158));
  inv1   g1086(.a(n1158), .O(n1159));
  nor2   g1087(.a(n740), .b(n272), .O(n1160));
  nor2   g1088(.a(n732), .b(n767), .O(n1161));
  nor2   g1089(.a(n1161), .b(n1160), .O(n1162));
  inv1   g1090(.a(n1162), .O(n1163));
  nor2   g1091(.a(n722), .b(n761), .O(n1164));
  nor2   g1092(.a(n727), .b(n320), .O(n1165));
  nor2   g1093(.a(n1165), .b(n1164), .O(n1166));
  inv1   g1094(.a(n1166), .O(n1167));
  nor2   g1095(.a(n1167), .b(n1163), .O(n1168));
  inv1   g1096(.a(n1168), .O(n1169));
  nor2   g1097(.a(n1169), .b(n1159), .O(n1170));
  inv1   g1098(.a(n1170), .O(n1171));
  nor2   g1099(.a(n1171), .b(n1157), .O(n1172));
  nor2   g1100(.a(n1172), .b(n1150), .O(n1173));
  nor2   g1101(.a(n1173), .b(n695), .O(n1174));
  nor2   g1102(.a(n675), .b(n180), .O(n1175));
  nor2   g1103(.a(n133), .b(G97), .O(n1176));
  nor2   g1104(.a(n1176), .b(n681), .O(n1177));
  inv1   g1105(.a(n1177), .O(n1178));
  nor2   g1106(.a(n1178), .b(n1175), .O(n1179));
  nor2   g1107(.a(n1179), .b(n672), .O(n1180));
  nor2   g1108(.a(n1180), .b(n694), .O(n1181));
  inv1   g1109(.a(n1181), .O(n1182));
  nor2   g1110(.a(n1182), .b(n1174), .O(n1183));
  inv1   g1111(.a(n1183), .O(n1184));
  nor2   g1112(.a(n1184), .b(n1128), .O(n1185));
  nor2   g1113(.a(n1185), .b(n1127), .O(n1186));
  inv1   g1114(.a(n1186), .O(n1187));
  nor2   g1115(.a(n1187), .b(n1126), .O(n1188));
  inv1   g1116(.a(n1188), .O(G390));
  nor2   g1117(.a(n796), .b(n857), .O(n1190));
  inv1   g1118(.a(n1190), .O(n1191));
  nor2   g1119(.a(n1191), .b(n879), .O(n1192));
  inv1   g1120(.a(n881), .O(n1193));
  inv1   g1121(.a(n886), .O(n1194));
  nor2   g1122(.a(n1194), .b(n1193), .O(n1195));
  nor2   g1123(.a(n1195), .b(n887), .O(n1196));
  inv1   g1124(.a(n1196), .O(n1197));
  nor2   g1125(.a(n1197), .b(n1192), .O(n1198));
  inv1   g1126(.a(n1192), .O(n1199));
  nor2   g1127(.a(n1196), .b(n1199), .O(n1200));
  nor2   g1128(.a(n1200), .b(n1198), .O(n1201));
  inv1   g1129(.a(n1201), .O(n1202));
  nor2   g1130(.a(n648), .b(n575), .O(n1203));
  nor2   g1131(.a(n1203), .b(n596), .O(n1204));
  inv1   g1132(.a(n1204), .O(n1205));
  inv1   g1133(.a(n874), .O(n1206));
  inv1   g1134(.a(n879), .O(n1207));
  nor2   g1135(.a(n1190), .b(n1207), .O(n1208));
  nor2   g1136(.a(n1208), .b(n1192), .O(n1209));
  inv1   g1137(.a(n1209), .O(n1210));
  nor2   g1138(.a(n1210), .b(n1206), .O(n1211));
  nor2   g1139(.a(n1209), .b(n874), .O(n1212));
  nor2   g1140(.a(n1212), .b(n1211), .O(n1213));
  nor2   g1141(.a(n1213), .b(n1205), .O(n1214));
  nor2   g1142(.a(n1214), .b(n1202), .O(n1215));
  inv1   g1143(.a(n1214), .O(n1216));
  nor2   g1144(.a(n1216), .b(n1201), .O(n1217));
  nor2   g1145(.a(n1217), .b(n657), .O(n1218));
  inv1   g1146(.a(n1218), .O(n1219));
  nor2   g1147(.a(n1219), .b(n1215), .O(n1220));
  nor2   g1148(.a(n1201), .b(n691), .O(n1221));
  nor2   g1149(.a(n1194), .b(n791), .O(n1222));
  nor2   g1150(.a(n702), .b(n106), .O(n1223));
  nor2   g1151(.a(n708), .b(n453), .O(n1224));
  inv1   g1152(.a(G125), .O(n1225));
  nor2   g1153(.a(n712), .b(n1225), .O(n1226));
  nor2   g1154(.a(n1226), .b(n1224), .O(n1227));
  inv1   g1155(.a(n1227), .O(n1228));
  nor2   g1156(.a(n1228), .b(n1223), .O(n1229));
  inv1   g1157(.a(n1229), .O(n1230));
  inv1   g1158(.a(G128), .O(n1231));
  nor2   g1159(.a(n722), .b(n1231), .O(n1232));
  nor2   g1160(.a(n1232), .b(G33), .O(n1233));
  inv1   g1161(.a(n1233), .O(n1234));
  nor2   g1162(.a(n727), .b(n807), .O(n1235));
  nor2   g1163(.a(n732), .b(n801), .O(n1236));
  nor2   g1164(.a(n1236), .b(n1235), .O(n1237));
  inv1   g1165(.a(n1237), .O(n1238));
  nor2   g1166(.a(n737), .b(n812), .O(n1239));
  nor2   g1167(.a(n740), .b(n404), .O(n1240));
  nor2   g1168(.a(n1240), .b(n1239), .O(n1241));
  inv1   g1169(.a(n1241), .O(n1242));
  nor2   g1170(.a(n1242), .b(n1238), .O(n1243));
  inv1   g1171(.a(n1243), .O(n1244));
  nor2   g1172(.a(n1244), .b(n1234), .O(n1245));
  inv1   g1173(.a(n1245), .O(n1246));
  nor2   g1174(.a(n1246), .b(n1230), .O(n1247));
  nor2   g1175(.a(n732), .b(n88), .O(n1248));
  nor2   g1176(.a(n712), .b(n375), .O(n1249));
  nor2   g1177(.a(n722), .b(n272), .O(n1250));
  nor2   g1178(.a(n1250), .b(n1249), .O(n1251));
  inv1   g1179(.a(n1251), .O(n1252));
  nor2   g1180(.a(n1252), .b(n1248), .O(n1253));
  inv1   g1181(.a(n1253), .O(n1254));
  nor2   g1182(.a(n741), .b(n197), .O(n1255));
  inv1   g1183(.a(n1255), .O(n1256));
  nor2   g1184(.a(n1129), .b(n799), .O(n1257));
  inv1   g1185(.a(n1257), .O(n1258));
  nor2   g1186(.a(n737), .b(n96), .O(n1259));
  nor2   g1187(.a(n727), .b(n103), .O(n1260));
  nor2   g1188(.a(n1260), .b(n1259), .O(n1261));
  inv1   g1189(.a(n1261), .O(n1262));
  nor2   g1190(.a(n1262), .b(n1258), .O(n1263));
  inv1   g1191(.a(n1263), .O(n1264));
  nor2   g1192(.a(n1264), .b(n1256), .O(n1265));
  inv1   g1193(.a(n1265), .O(n1266));
  nor2   g1194(.a(n1266), .b(n1254), .O(n1267));
  nor2   g1195(.a(n1267), .b(n1247), .O(n1268));
  nor2   g1196(.a(n1268), .b(n695), .O(n1269));
  nor2   g1197(.a(n850), .b(G58), .O(n1270));
  nor2   g1198(.a(n1270), .b(n694), .O(n1271));
  inv1   g1199(.a(n1271), .O(n1272));
  nor2   g1200(.a(n1272), .b(n1269), .O(n1273));
  inv1   g1201(.a(n1273), .O(n1274));
  nor2   g1202(.a(n1274), .b(n1222), .O(n1275));
  nor2   g1203(.a(n1275), .b(n1221), .O(n1276));
  inv1   g1204(.a(n1276), .O(n1277));
  nor2   g1205(.a(n1277), .b(n1220), .O(n1278));
  inv1   g1206(.a(n1278), .O(G378));
  nor2   g1207(.a(n1217), .b(n1205), .O(n1280));
  inv1   g1208(.a(n895), .O(n1281));
  nor2   g1209(.a(n1281), .b(n619), .O(n1282));
  nor2   g1210(.a(n1282), .b(n901), .O(n1283));
  inv1   g1211(.a(n1282), .O(n1284));
  nor2   g1212(.a(n1284), .b(n888), .O(n1285));
  nor2   g1213(.a(n1285), .b(n1283), .O(n1286));
  inv1   g1214(.a(n1286), .O(n1287));
  nor2   g1215(.a(n605), .b(n419), .O(n1288));
  nor2   g1216(.a(n1288), .b(n452), .O(n1289));
  inv1   g1217(.a(n444), .O(n1290));
  inv1   g1218(.a(n1288), .O(n1291));
  nor2   g1219(.a(n1291), .b(n1290), .O(n1292));
  nor2   g1220(.a(n1292), .b(n1289), .O(n1293));
  inv1   g1221(.a(n1293), .O(n1294));
  nor2   g1222(.a(n1294), .b(n1287), .O(n1295));
  nor2   g1223(.a(n1293), .b(n1286), .O(n1296));
  nor2   g1224(.a(n1296), .b(n1295), .O(n1297));
  nor2   g1225(.a(n1297), .b(n657), .O(n1298));
  inv1   g1226(.a(n1298), .O(n1299));
  nor2   g1227(.a(n1299), .b(n1280), .O(n1300));
  nor2   g1228(.a(n1297), .b(n691), .O(n1301));
  nor2   g1229(.a(n1294), .b(n791), .O(n1302));
  nor2   g1230(.a(n702), .b(n453), .O(n1303));
  inv1   g1231(.a(G124), .O(n1304));
  nor2   g1232(.a(n712), .b(n1304), .O(n1305));
  nor2   g1233(.a(n708), .b(n404), .O(n1306));
  nor2   g1234(.a(n1306), .b(n1305), .O(n1307));
  inv1   g1235(.a(n1307), .O(n1308));
  nor2   g1236(.a(n1308), .b(n1303), .O(n1309));
  inv1   g1237(.a(n1309), .O(n1310));
  nor2   g1238(.a(n722), .b(n1225), .O(n1311));
  nor2   g1239(.a(G41), .b(G33), .O(n1312));
  inv1   g1240(.a(n1312), .O(n1313));
  nor2   g1241(.a(n1313), .b(n1311), .O(n1314));
  inv1   g1242(.a(n1314), .O(n1315));
  nor2   g1243(.a(n727), .b(n801), .O(n1316));
  nor2   g1244(.a(n732), .b(n1231), .O(n1317));
  nor2   g1245(.a(n1317), .b(n1316), .O(n1318));
  inv1   g1246(.a(n1318), .O(n1319));
  nor2   g1247(.a(n737), .b(n807), .O(n1320));
  nor2   g1248(.a(n740), .b(n812), .O(n1321));
  nor2   g1249(.a(n1321), .b(n1320), .O(n1322));
  inv1   g1250(.a(n1322), .O(n1323));
  nor2   g1251(.a(n1323), .b(n1319), .O(n1324));
  inv1   g1252(.a(n1324), .O(n1325));
  nor2   g1253(.a(n1325), .b(n1315), .O(n1326));
  inv1   g1254(.a(n1326), .O(n1327));
  nor2   g1255(.a(n1327), .b(n1310), .O(n1328));
  nor2   g1256(.a(G50), .b(n198), .O(n1329));
  nor2   g1257(.a(n727), .b(n96), .O(n1330));
  nor2   g1258(.a(n732), .b(n103), .O(n1331));
  nor2   g1259(.a(n712), .b(n272), .O(n1332));
  nor2   g1260(.a(n1332), .b(n1331), .O(n1333));
  inv1   g1261(.a(n1333), .O(n1334));
  nor2   g1262(.a(n1334), .b(n1330), .O(n1335));
  inv1   g1263(.a(n1335), .O(n1336));
  nor2   g1264(.a(G41), .b(n197), .O(n1337));
  inv1   g1265(.a(n1337), .O(n1338));
  nor2   g1266(.a(n1338), .b(n980), .O(n1339));
  inv1   g1267(.a(n1339), .O(n1340));
  nor2   g1268(.a(n702), .b(n93), .O(n1341));
  nor2   g1269(.a(n1341), .b(n1075), .O(n1342));
  inv1   g1270(.a(n1342), .O(n1343));
  nor2   g1271(.a(n722), .b(n88), .O(n1344));
  nor2   g1272(.a(n737), .b(n78), .O(n1345));
  nor2   g1273(.a(n1345), .b(n1344), .O(n1346));
  inv1   g1274(.a(n1346), .O(n1347));
  nor2   g1275(.a(n1347), .b(n1343), .O(n1348));
  inv1   g1276(.a(n1348), .O(n1349));
  nor2   g1277(.a(n1349), .b(n1340), .O(n1350));
  inv1   g1278(.a(n1350), .O(n1351));
  nor2   g1279(.a(n1351), .b(n1336), .O(n1352));
  nor2   g1280(.a(n1352), .b(n1329), .O(n1353));
  inv1   g1281(.a(n1353), .O(n1354));
  nor2   g1282(.a(n1354), .b(n1328), .O(n1355));
  nor2   g1283(.a(n1355), .b(n695), .O(n1356));
  nor2   g1284(.a(n850), .b(G50), .O(n1357));
  nor2   g1285(.a(n1357), .b(n694), .O(n1358));
  inv1   g1286(.a(n1358), .O(n1359));
  nor2   g1287(.a(n1359), .b(n1356), .O(n1360));
  inv1   g1288(.a(n1360), .O(n1361));
  nor2   g1289(.a(n1361), .b(n1302), .O(n1362));
  nor2   g1290(.a(n1362), .b(n1301), .O(n1363));
  inv1   g1291(.a(n1363), .O(n1364));
  nor2   g1292(.a(n1364), .b(n1300), .O(n1365));
  inv1   g1293(.a(n1365), .O(G375));
  inv1   g1294(.a(n1213), .O(n1367));
  nor2   g1295(.a(n1367), .b(n1204), .O(n1368));
  nor2   g1296(.a(n1214), .b(n657), .O(n1369));
  inv1   g1297(.a(n1369), .O(n1370));
  nor2   g1298(.a(n1370), .b(n1368), .O(n1371));
  nor2   g1299(.a(n1213), .b(n691), .O(n1372));
  nor2   g1300(.a(n1207), .b(n791), .O(n1373));
  nor2   g1301(.a(n708), .b(n106), .O(n1374));
  nor2   g1302(.a(n712), .b(n1231), .O(n1375));
  nor2   g1303(.a(n737), .b(n404), .O(n1376));
  nor2   g1304(.a(n1376), .b(n1375), .O(n1377));
  inv1   g1305(.a(n1377), .O(n1378));
  nor2   g1306(.a(n1378), .b(n1374), .O(n1379));
  inv1   g1307(.a(n1379), .O(n1380));
  nor2   g1308(.a(n1341), .b(G33), .O(n1381));
  inv1   g1309(.a(n1381), .O(n1382));
  nor2   g1310(.a(n740), .b(n453), .O(n1383));
  nor2   g1311(.a(n732), .b(n807), .O(n1384));
  nor2   g1312(.a(n1384), .b(n1383), .O(n1385));
  inv1   g1313(.a(n1385), .O(n1386));
  nor2   g1314(.a(n722), .b(n801), .O(n1387));
  nor2   g1315(.a(n727), .b(n812), .O(n1388));
  nor2   g1316(.a(n1388), .b(n1387), .O(n1389));
  inv1   g1317(.a(n1389), .O(n1390));
  nor2   g1318(.a(n1390), .b(n1386), .O(n1391));
  inv1   g1319(.a(n1391), .O(n1392));
  nor2   g1320(.a(n1392), .b(n1382), .O(n1393));
  inv1   g1321(.a(n1393), .O(n1394));
  nor2   g1322(.a(n1394), .b(n1380), .O(n1395));
  nor2   g1323(.a(n727), .b(n88), .O(n1396));
  nor2   g1324(.a(n732), .b(n272), .O(n1397));
  nor2   g1325(.a(n740), .b(n96), .O(n1398));
  nor2   g1326(.a(n1398), .b(n1397), .O(n1399));
  inv1   g1327(.a(n1399), .O(n1400));
  nor2   g1328(.a(n1400), .b(n1396), .O(n1401));
  inv1   g1329(.a(n1401), .O(n1402));
  nor2   g1330(.a(n979), .b(n197), .O(n1403));
  inv1   g1331(.a(n1403), .O(n1404));
  nor2   g1332(.a(n712), .b(n320), .O(n1405));
  nor2   g1333(.a(n1405), .b(n1066), .O(n1406));
  inv1   g1334(.a(n1406), .O(n1407));
  nor2   g1335(.a(n722), .b(n375), .O(n1408));
  nor2   g1336(.a(n737), .b(n103), .O(n1409));
  nor2   g1337(.a(n1409), .b(n1408), .O(n1410));
  inv1   g1338(.a(n1410), .O(n1411));
  nor2   g1339(.a(n1411), .b(n1407), .O(n1412));
  inv1   g1340(.a(n1412), .O(n1413));
  nor2   g1341(.a(n1413), .b(n1404), .O(n1414));
  inv1   g1342(.a(n1414), .O(n1415));
  nor2   g1343(.a(n1415), .b(n1402), .O(n1416));
  nor2   g1344(.a(n1416), .b(n1395), .O(n1417));
  nor2   g1345(.a(n1417), .b(n695), .O(n1418));
  nor2   g1346(.a(n850), .b(G68), .O(n1419));
  nor2   g1347(.a(n1419), .b(n694), .O(n1420));
  inv1   g1348(.a(n1420), .O(n1421));
  nor2   g1349(.a(n1421), .b(n1418), .O(n1422));
  inv1   g1350(.a(n1422), .O(n1423));
  nor2   g1351(.a(n1423), .b(n1373), .O(n1424));
  nor2   g1352(.a(n1424), .b(n1372), .O(n1425));
  inv1   g1353(.a(n1425), .O(n1426));
  nor2   g1354(.a(n1426), .b(n1371), .O(n1427));
  inv1   g1355(.a(n1427), .O(G381));
  nor2   g1356(.a(G384), .b(G396), .O(n1429));
  inv1   g1357(.a(n1429), .O(n1430));
  nor2   g1358(.a(n1430), .b(G393), .O(n1431));
  inv1   g1359(.a(n1431), .O(n1432));
  nor2   g1360(.a(n1432), .b(G390), .O(n1433));
  inv1   g1361(.a(n1433), .O(n1434));
  nor2   g1362(.a(n1434), .b(G387), .O(n1435));
  inv1   g1363(.a(n1435), .O(n1436));
  nor2   g1364(.a(n1436), .b(G381), .O(n1437));
  inv1   g1365(.a(n1437), .O(n1438));
  nor2   g1366(.a(n1438), .b(G378), .O(n1439));
  inv1   g1367(.a(n1439), .O(n1440));
  nor2   g1368(.a(n1440), .b(G375), .O(n1441));
  inv1   g1369(.a(n1441), .O(G407));
  nor2   g1370(.a(G343), .b(n601), .O(n1443));
  inv1   g1371(.a(n1443), .O(n1444));
  nor2   g1372(.a(n1444), .b(G378), .O(n1445));
  inv1   g1373(.a(n1445), .O(n1446));
  nor2   g1374(.a(n1446), .b(G375), .O(n1447));
  nor2   g1375(.a(n1441), .b(n601), .O(n1448));
  inv1   g1376(.a(n1448), .O(n1449));
  nor2   g1377(.a(n1449), .b(n1447), .O(n1450));
  inv1   g1378(.a(n1450), .O(G409));
  nor2   g1379(.a(n1365), .b(G378), .O(n1452));
  nor2   g1380(.a(G375), .b(n1278), .O(n1453));
  nor2   g1381(.a(n1453), .b(n1452), .O(n1454));
  inv1   g1382(.a(n1454), .O(n1455));
  nor2   g1383(.a(n1455), .b(n1443), .O(n1456));
  nor2   g1384(.a(n1444), .b(G2897), .O(n1457));
  nor2   g1385(.a(n1457), .b(n1456), .O(n1458));
  nor2   g1386(.a(G390), .b(n1040), .O(n1459));
  nor2   g1387(.a(n1188), .b(G387), .O(n1460));
  nor2   g1388(.a(n1460), .b(n1459), .O(n1461));
  inv1   g1389(.a(n1461), .O(n1462));
  nor2   g1390(.a(n1462), .b(n1120), .O(n1463));
  nor2   g1391(.a(n1461), .b(G393), .O(n1464));
  nor2   g1392(.a(n1464), .b(n1463), .O(n1465));
  inv1   g1393(.a(n1465), .O(n1466));
  nor2   g1394(.a(n1427), .b(G384), .O(n1467));
  nor2   g1395(.a(G381), .b(n868), .O(n1468));
  nor2   g1396(.a(n1468), .b(n1467), .O(n1469));
  inv1   g1397(.a(n1469), .O(n1470));
  nor2   g1398(.a(n1470), .b(n788), .O(n1471));
  nor2   g1399(.a(n1469), .b(G396), .O(n1472));
  nor2   g1400(.a(n1472), .b(n1471), .O(n1473));
  inv1   g1401(.a(n1473), .O(n1474));
  nor2   g1402(.a(n1474), .b(n1466), .O(n1475));
  nor2   g1403(.a(n1473), .b(n1465), .O(n1476));
  nor2   g1404(.a(n1476), .b(n1475), .O(n1477));
  inv1   g1405(.a(n1477), .O(n1478));
  nor2   g1406(.a(n1478), .b(n1458), .O(n1479));
  inv1   g1407(.a(n1458), .O(n1480));
  nor2   g1408(.a(n1477), .b(n1480), .O(n1481));
  nor2   g1409(.a(n1481), .b(n1479), .O(G405));
  nor2   g1410(.a(n1478), .b(n1455), .O(n1483));
  nor2   g1411(.a(n1477), .b(n1454), .O(n1484));
  nor2   g1412(.a(n1484), .b(n1483), .O(G402));
endmodule


