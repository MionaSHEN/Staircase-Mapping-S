// Benchmark "c1355_blif" written by ABC on Sun Apr 14 20:05:53 2019

module c1355_blif  ( 
    G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat,
    G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat,
    G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat,
    G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat,
    G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat,
    G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat,
    G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat,
    G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat,
    G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat,
    G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n446, n447, n448, n449, n450,
    n452, n453, n454, n455, n456, n458, n459, n460, n461, n462, n464, n465,
    n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n477, n478,
    n479, n480, n481, n483, n484, n485, n486, n487, n489, n490, n491, n492,
    n493, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
    n506, n508, n509, n510, n511, n512, n514, n515, n516, n517, n518, n520,
    n521, n522, n523, n524, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n538, n539, n540, n541, n542, n544, n545, n546, n547,
    n548, n550, n551, n552, n553, n554, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
    n575, n576, n577, n578, n579, n581, n582, n583, n584, n585, n587, n588,
    n589, n590, n591, n593, n594, n595, n596, n597, n598, n599, n600, n601,
    n602, n604, n605, n606, n607, n608, n610, n611, n612, n613, n614, n616,
    n617, n618, n619, n620, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n632, n633, n634, n635, n636, n638, n639, n640, n641, n642, n644,
    n645, n646, n647, n648, n650, n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n661, n662, n663, n664, n665, n667, n668, n669, n670, n671,
    n673, n674, n675, n676, n677;
  inv1   g000(.a(G1gat), .O(n74));
  inv1   g001(.a(G113gat), .O(n75));
  nor2   g002(.a(G134gat), .b(n75), .O(n76));
  inv1   g003(.a(G134gat), .O(n77));
  nor2   g004(.a(n77), .b(G113gat), .O(n78));
  nor2   g005(.a(n78), .b(n76), .O(n79));
  inv1   g006(.a(n79), .O(n80));
  inv1   g007(.a(G120gat), .O(n81));
  nor2   g008(.a(G127gat), .b(n81), .O(n82));
  inv1   g009(.a(G127gat), .O(n83));
  nor2   g010(.a(n83), .b(G120gat), .O(n84));
  nor2   g011(.a(n84), .b(n82), .O(n85));
  nor2   g012(.a(n85), .b(n80), .O(n86));
  inv1   g013(.a(n85), .O(n87));
  nor2   g014(.a(n87), .b(n79), .O(n88));
  nor2   g015(.a(n88), .b(n86), .O(n89));
  inv1   g016(.a(n89), .O(n90));
  inv1   g017(.a(G225gat), .O(n91));
  inv1   g018(.a(G233gat), .O(n92));
  nor2   g019(.a(n92), .b(n91), .O(n93));
  inv1   g020(.a(n93), .O(n94));
  nor2   g021(.a(n94), .b(n90), .O(n95));
  nor2   g022(.a(n93), .b(n89), .O(n96));
  nor2   g023(.a(n96), .b(n95), .O(n97));
  inv1   g024(.a(n97), .O(n98));
  inv1   g025(.a(G141gat), .O(n99));
  nor2   g026(.a(G162gat), .b(n99), .O(n100));
  inv1   g027(.a(G162gat), .O(n101));
  nor2   g028(.a(n101), .b(G141gat), .O(n102));
  nor2   g029(.a(n102), .b(n100), .O(n103));
  inv1   g030(.a(n103), .O(n104));
  inv1   g031(.a(G148gat), .O(n105));
  nor2   g032(.a(G155gat), .b(n105), .O(n106));
  inv1   g033(.a(G155gat), .O(n107));
  nor2   g034(.a(n107), .b(G148gat), .O(n108));
  nor2   g035(.a(n108), .b(n106), .O(n109));
  nor2   g036(.a(n109), .b(n104), .O(n110));
  inv1   g037(.a(n109), .O(n111));
  nor2   g038(.a(n111), .b(n103), .O(n112));
  nor2   g039(.a(n112), .b(n110), .O(n113));
  nor2   g040(.a(G85gat), .b(n74), .O(n114));
  inv1   g041(.a(G85gat), .O(n115));
  nor2   g042(.a(n115), .b(G1gat), .O(n116));
  nor2   g043(.a(n116), .b(n114), .O(n117));
  inv1   g044(.a(n117), .O(n118));
  inv1   g045(.a(G29gat), .O(n119));
  nor2   g046(.a(G57gat), .b(n119), .O(n120));
  inv1   g047(.a(G57gat), .O(n121));
  nor2   g048(.a(n121), .b(G29gat), .O(n122));
  nor2   g049(.a(n122), .b(n120), .O(n123));
  nor2   g050(.a(n123), .b(n118), .O(n124));
  inv1   g051(.a(n123), .O(n125));
  nor2   g052(.a(n125), .b(n117), .O(n126));
  nor2   g053(.a(n126), .b(n124), .O(n127));
  inv1   g054(.a(n127), .O(n128));
  nor2   g055(.a(n128), .b(n113), .O(n129));
  inv1   g056(.a(n113), .O(n130));
  nor2   g057(.a(n127), .b(n130), .O(n131));
  nor2   g058(.a(n131), .b(n129), .O(n132));
  inv1   g059(.a(n132), .O(n133));
  nor2   g060(.a(n133), .b(n98), .O(n134));
  nor2   g061(.a(n132), .b(n97), .O(n135));
  nor2   g062(.a(n135), .b(n134), .O(n136));
  inv1   g063(.a(n136), .O(n137));
  inv1   g064(.a(G106gat), .O(n138));
  inv1   g065(.a(G78gat), .O(n139));
  inv1   g066(.a(G197gat), .O(n140));
  nor2   g067(.a(G218gat), .b(n140), .O(n141));
  inv1   g068(.a(G218gat), .O(n142));
  nor2   g069(.a(n142), .b(G197gat), .O(n143));
  nor2   g070(.a(n143), .b(n141), .O(n144));
  inv1   g071(.a(n144), .O(n145));
  inv1   g072(.a(G204gat), .O(n146));
  nor2   g073(.a(G211gat), .b(n146), .O(n147));
  inv1   g074(.a(G211gat), .O(n148));
  nor2   g075(.a(n148), .b(G204gat), .O(n149));
  nor2   g076(.a(n149), .b(n147), .O(n150));
  nor2   g077(.a(n150), .b(n145), .O(n151));
  inv1   g078(.a(n150), .O(n152));
  nor2   g079(.a(n152), .b(n144), .O(n153));
  nor2   g080(.a(n153), .b(n151), .O(n154));
  nor2   g081(.a(n154), .b(n139), .O(n155));
  inv1   g082(.a(n154), .O(n156));
  nor2   g083(.a(n156), .b(G78gat), .O(n157));
  nor2   g084(.a(n157), .b(n155), .O(n158));
  inv1   g085(.a(n158), .O(n159));
  nor2   g086(.a(n159), .b(n138), .O(n160));
  nor2   g087(.a(n158), .b(G106gat), .O(n161));
  nor2   g088(.a(n161), .b(n160), .O(n162));
  inv1   g089(.a(n162), .O(n163));
  inv1   g090(.a(G228gat), .O(n164));
  nor2   g091(.a(n92), .b(n164), .O(n165));
  inv1   g092(.a(n165), .O(n166));
  inv1   g093(.a(G22gat), .O(n167));
  nor2   g094(.a(G50gat), .b(n167), .O(n168));
  inv1   g095(.a(G50gat), .O(n169));
  nor2   g096(.a(n169), .b(G22gat), .O(n170));
  nor2   g097(.a(n170), .b(n168), .O(n171));
  nor2   g098(.a(n171), .b(n166), .O(n172));
  inv1   g099(.a(n171), .O(n173));
  nor2   g100(.a(n173), .b(n165), .O(n174));
  nor2   g101(.a(n174), .b(n172), .O(n175));
  nor2   g102(.a(n175), .b(n130), .O(n176));
  inv1   g103(.a(n175), .O(n177));
  nor2   g104(.a(n177), .b(n113), .O(n178));
  nor2   g105(.a(n178), .b(n176), .O(n179));
  inv1   g106(.a(n179), .O(n180));
  nor2   g107(.a(n180), .b(n163), .O(n181));
  nor2   g108(.a(n179), .b(n162), .O(n182));
  nor2   g109(.a(n182), .b(n181), .O(n183));
  inv1   g110(.a(n183), .O(n184));
  inv1   g111(.a(G99gat), .O(n185));
  inv1   g112(.a(G71gat), .O(n186));
  inv1   g113(.a(G169gat), .O(n187));
  nor2   g114(.a(G190gat), .b(n187), .O(n188));
  inv1   g115(.a(G190gat), .O(n189));
  nor2   g116(.a(n189), .b(G169gat), .O(n190));
  nor2   g117(.a(n190), .b(n188), .O(n191));
  inv1   g118(.a(n191), .O(n192));
  inv1   g119(.a(G176gat), .O(n193));
  nor2   g120(.a(G183gat), .b(n193), .O(n194));
  inv1   g121(.a(G183gat), .O(n195));
  nor2   g122(.a(n195), .b(G176gat), .O(n196));
  nor2   g123(.a(n196), .b(n194), .O(n197));
  nor2   g124(.a(n197), .b(n192), .O(n198));
  inv1   g125(.a(n197), .O(n199));
  nor2   g126(.a(n199), .b(n191), .O(n200));
  nor2   g127(.a(n200), .b(n198), .O(n201));
  nor2   g128(.a(n201), .b(n186), .O(n202));
  inv1   g129(.a(n201), .O(n203));
  nor2   g130(.a(n203), .b(G71gat), .O(n204));
  nor2   g131(.a(n204), .b(n202), .O(n205));
  inv1   g132(.a(n205), .O(n206));
  nor2   g133(.a(n206), .b(n185), .O(n207));
  nor2   g134(.a(n205), .b(G99gat), .O(n208));
  nor2   g135(.a(n208), .b(n207), .O(n209));
  inv1   g136(.a(n209), .O(n210));
  inv1   g137(.a(G227gat), .O(n211));
  nor2   g138(.a(n92), .b(n211), .O(n212));
  inv1   g139(.a(n212), .O(n213));
  inv1   g140(.a(G15gat), .O(n214));
  nor2   g141(.a(G43gat), .b(n214), .O(n215));
  inv1   g142(.a(G43gat), .O(n216));
  nor2   g143(.a(n216), .b(G15gat), .O(n217));
  nor2   g144(.a(n217), .b(n215), .O(n218));
  nor2   g145(.a(n218), .b(n213), .O(n219));
  inv1   g146(.a(n218), .O(n220));
  nor2   g147(.a(n220), .b(n212), .O(n221));
  nor2   g148(.a(n221), .b(n219), .O(n222));
  nor2   g149(.a(n222), .b(n90), .O(n223));
  inv1   g150(.a(n222), .O(n224));
  nor2   g151(.a(n224), .b(n89), .O(n225));
  nor2   g152(.a(n225), .b(n223), .O(n226));
  inv1   g153(.a(n226), .O(n227));
  nor2   g154(.a(n227), .b(n210), .O(n228));
  nor2   g155(.a(n226), .b(n209), .O(n229));
  nor2   g156(.a(n229), .b(n228), .O(n230));
  nor2   g157(.a(n230), .b(n184), .O(n231));
  inv1   g158(.a(n230), .O(n232));
  nor2   g159(.a(n232), .b(n183), .O(n233));
  nor2   g160(.a(n233), .b(n231), .O(n234));
  inv1   g161(.a(G226gat), .O(n235));
  nor2   g162(.a(n92), .b(n235), .O(n236));
  inv1   g163(.a(n236), .O(n237));
  nor2   g164(.a(n237), .b(n156), .O(n238));
  nor2   g165(.a(n236), .b(n154), .O(n239));
  nor2   g166(.a(n239), .b(n238), .O(n240));
  inv1   g167(.a(n240), .O(n241));
  inv1   g168(.a(G64gat), .O(n242));
  nor2   g169(.a(G92gat), .b(n242), .O(n243));
  inv1   g170(.a(G92gat), .O(n244));
  nor2   g171(.a(n244), .b(G64gat), .O(n245));
  nor2   g172(.a(n245), .b(n243), .O(n246));
  inv1   g173(.a(n246), .O(n247));
  inv1   g174(.a(G8gat), .O(n248));
  nor2   g175(.a(G36gat), .b(n248), .O(n249));
  inv1   g176(.a(G36gat), .O(n250));
  nor2   g177(.a(n250), .b(G8gat), .O(n251));
  nor2   g178(.a(n251), .b(n249), .O(n252));
  nor2   g179(.a(n252), .b(n247), .O(n253));
  inv1   g180(.a(n252), .O(n254));
  nor2   g181(.a(n254), .b(n246), .O(n255));
  nor2   g182(.a(n255), .b(n253), .O(n256));
  nor2   g183(.a(n256), .b(n203), .O(n257));
  inv1   g184(.a(n256), .O(n258));
  nor2   g185(.a(n258), .b(n201), .O(n259));
  nor2   g186(.a(n259), .b(n257), .O(n260));
  inv1   g187(.a(n260), .O(n261));
  nor2   g188(.a(n261), .b(n241), .O(n262));
  nor2   g189(.a(n260), .b(n240), .O(n263));
  nor2   g190(.a(n263), .b(n262), .O(n264));
  nor2   g191(.a(n264), .b(n136), .O(n265));
  inv1   g192(.a(n265), .O(n266));
  nor2   g193(.a(n266), .b(n234), .O(n267));
  inv1   g194(.a(n264), .O(n268));
  nor2   g195(.a(n268), .b(n136), .O(n269));
  inv1   g196(.a(n269), .O(n270));
  nor2   g197(.a(n270), .b(n230), .O(n271));
  nor2   g198(.a(n264), .b(n137), .O(n272));
  inv1   g199(.a(n272), .O(n273));
  nor2   g200(.a(n273), .b(n230), .O(n274));
  nor2   g201(.a(n274), .b(n271), .O(n275));
  nor2   g202(.a(n275), .b(n183), .O(n276));
  nor2   g203(.a(n276), .b(n267), .O(n277));
  inv1   g204(.a(G229gat), .O(n278));
  nor2   g205(.a(n92), .b(n278), .O(n279));
  inv1   g206(.a(n279), .O(n280));
  nor2   g207(.a(G50gat), .b(n119), .O(n281));
  nor2   g208(.a(n169), .b(G29gat), .O(n282));
  nor2   g209(.a(n282), .b(n281), .O(n283));
  inv1   g210(.a(n283), .O(n284));
  nor2   g211(.a(G43gat), .b(n250), .O(n285));
  nor2   g212(.a(n216), .b(G36gat), .O(n286));
  nor2   g213(.a(n286), .b(n285), .O(n287));
  nor2   g214(.a(n287), .b(n284), .O(n288));
  inv1   g215(.a(n287), .O(n289));
  nor2   g216(.a(n289), .b(n283), .O(n290));
  nor2   g217(.a(n290), .b(n288), .O(n291));
  inv1   g218(.a(n291), .O(n292));
  nor2   g219(.a(n292), .b(n280), .O(n293));
  nor2   g220(.a(n291), .b(n279), .O(n294));
  nor2   g221(.a(n294), .b(n293), .O(n295));
  inv1   g222(.a(n295), .O(n296));
  nor2   g223(.a(G22gat), .b(n74), .O(n297));
  nor2   g224(.a(n167), .b(G1gat), .O(n298));
  nor2   g225(.a(n298), .b(n297), .O(n299));
  inv1   g226(.a(n299), .O(n300));
  nor2   g227(.a(G15gat), .b(n248), .O(n301));
  nor2   g228(.a(n214), .b(G8gat), .O(n302));
  nor2   g229(.a(n302), .b(n301), .O(n303));
  nor2   g230(.a(n303), .b(n300), .O(n304));
  inv1   g231(.a(n303), .O(n305));
  nor2   g232(.a(n305), .b(n299), .O(n306));
  nor2   g233(.a(n306), .b(n304), .O(n307));
  inv1   g234(.a(n307), .O(n308));
  nor2   g235(.a(G197gat), .b(n187), .O(n309));
  nor2   g236(.a(n140), .b(G169gat), .O(n310));
  nor2   g237(.a(n310), .b(n309), .O(n311));
  inv1   g238(.a(n311), .O(n312));
  nor2   g239(.a(G141gat), .b(n75), .O(n313));
  nor2   g240(.a(n99), .b(G113gat), .O(n314));
  nor2   g241(.a(n314), .b(n313), .O(n315));
  nor2   g242(.a(n315), .b(n312), .O(n316));
  inv1   g243(.a(n315), .O(n317));
  nor2   g244(.a(n317), .b(n311), .O(n318));
  nor2   g245(.a(n318), .b(n316), .O(n319));
  nor2   g246(.a(n319), .b(n308), .O(n320));
  inv1   g247(.a(n319), .O(n321));
  nor2   g248(.a(n321), .b(n307), .O(n322));
  nor2   g249(.a(n322), .b(n320), .O(n323));
  inv1   g250(.a(n323), .O(n324));
  nor2   g251(.a(n324), .b(n296), .O(n325));
  nor2   g252(.a(n323), .b(n295), .O(n326));
  nor2   g253(.a(n326), .b(n325), .O(n327));
  inv1   g254(.a(n327), .O(n328));
  inv1   g255(.a(G230gat), .O(n329));
  nor2   g256(.a(n92), .b(n329), .O(n330));
  inv1   g257(.a(n330), .O(n331));
  nor2   g258(.a(G106gat), .b(n115), .O(n332));
  nor2   g259(.a(n138), .b(G85gat), .O(n333));
  nor2   g260(.a(n333), .b(n332), .O(n334));
  inv1   g261(.a(n334), .O(n335));
  nor2   g262(.a(G99gat), .b(n244), .O(n336));
  nor2   g263(.a(n185), .b(G92gat), .O(n337));
  nor2   g264(.a(n337), .b(n336), .O(n338));
  nor2   g265(.a(n338), .b(n335), .O(n339));
  inv1   g266(.a(n338), .O(n340));
  nor2   g267(.a(n340), .b(n334), .O(n341));
  nor2   g268(.a(n341), .b(n339), .O(n342));
  inv1   g269(.a(n342), .O(n343));
  nor2   g270(.a(n343), .b(n331), .O(n344));
  nor2   g271(.a(n342), .b(n330), .O(n345));
  nor2   g272(.a(n345), .b(n344), .O(n346));
  inv1   g273(.a(n346), .O(n347));
  nor2   g274(.a(G78gat), .b(n121), .O(n348));
  nor2   g275(.a(n139), .b(G57gat), .O(n349));
  nor2   g276(.a(n349), .b(n348), .O(n350));
  inv1   g277(.a(n350), .O(n351));
  nor2   g278(.a(G71gat), .b(n242), .O(n352));
  nor2   g279(.a(n186), .b(G64gat), .O(n353));
  nor2   g280(.a(n353), .b(n352), .O(n354));
  nor2   g281(.a(n354), .b(n351), .O(n355));
  inv1   g282(.a(n354), .O(n356));
  nor2   g283(.a(n356), .b(n350), .O(n357));
  nor2   g284(.a(n357), .b(n355), .O(n358));
  inv1   g285(.a(n358), .O(n359));
  nor2   g286(.a(G204gat), .b(n193), .O(n360));
  nor2   g287(.a(n146), .b(G176gat), .O(n361));
  nor2   g288(.a(n361), .b(n360), .O(n362));
  inv1   g289(.a(n362), .O(n363));
  nor2   g290(.a(G148gat), .b(n81), .O(n364));
  nor2   g291(.a(n105), .b(G120gat), .O(n365));
  nor2   g292(.a(n365), .b(n364), .O(n366));
  nor2   g293(.a(n366), .b(n363), .O(n367));
  inv1   g294(.a(n366), .O(n368));
  nor2   g295(.a(n368), .b(n362), .O(n369));
  nor2   g296(.a(n369), .b(n367), .O(n370));
  nor2   g297(.a(n370), .b(n359), .O(n371));
  inv1   g298(.a(n370), .O(n372));
  nor2   g299(.a(n372), .b(n358), .O(n373));
  nor2   g300(.a(n373), .b(n371), .O(n374));
  inv1   g301(.a(n374), .O(n375));
  nor2   g302(.a(n375), .b(n347), .O(n376));
  nor2   g303(.a(n374), .b(n346), .O(n377));
  nor2   g304(.a(n377), .b(n376), .O(n378));
  nor2   g305(.a(n378), .b(n328), .O(n379));
  inv1   g306(.a(n379), .O(n380));
  nor2   g307(.a(n342), .b(n189), .O(n381));
  nor2   g308(.a(n343), .b(G190gat), .O(n382));
  nor2   g309(.a(n382), .b(n381), .O(n383));
  inv1   g310(.a(n383), .O(n384));
  nor2   g311(.a(n384), .b(n142), .O(n385));
  nor2   g312(.a(n383), .b(G218gat), .O(n386));
  nor2   g313(.a(n386), .b(n385), .O(n387));
  inv1   g314(.a(n387), .O(n388));
  inv1   g315(.a(G232gat), .O(n389));
  nor2   g316(.a(n92), .b(n389), .O(n390));
  inv1   g317(.a(n390), .O(n391));
  nor2   g318(.a(G162gat), .b(n77), .O(n392));
  nor2   g319(.a(n101), .b(G134gat), .O(n393));
  nor2   g320(.a(n393), .b(n392), .O(n394));
  nor2   g321(.a(n394), .b(n391), .O(n395));
  inv1   g322(.a(n394), .O(n396));
  nor2   g323(.a(n396), .b(n390), .O(n397));
  nor2   g324(.a(n397), .b(n395), .O(n398));
  nor2   g325(.a(n398), .b(n292), .O(n399));
  inv1   g326(.a(n398), .O(n400));
  nor2   g327(.a(n400), .b(n291), .O(n401));
  nor2   g328(.a(n401), .b(n399), .O(n402));
  inv1   g329(.a(n402), .O(n403));
  nor2   g330(.a(n403), .b(n388), .O(n404));
  nor2   g331(.a(n402), .b(n387), .O(n405));
  nor2   g332(.a(n405), .b(n404), .O(n406));
  nor2   g333(.a(n358), .b(n195), .O(n407));
  nor2   g334(.a(n359), .b(G183gat), .O(n408));
  nor2   g335(.a(n408), .b(n407), .O(n409));
  inv1   g336(.a(n409), .O(n410));
  nor2   g337(.a(n410), .b(n148), .O(n411));
  nor2   g338(.a(n409), .b(G211gat), .O(n412));
  nor2   g339(.a(n412), .b(n411), .O(n413));
  inv1   g340(.a(n413), .O(n414));
  inv1   g341(.a(G231gat), .O(n415));
  nor2   g342(.a(n92), .b(n415), .O(n416));
  inv1   g343(.a(n416), .O(n417));
  nor2   g344(.a(G155gat), .b(n83), .O(n418));
  nor2   g345(.a(n107), .b(G127gat), .O(n419));
  nor2   g346(.a(n419), .b(n418), .O(n420));
  nor2   g347(.a(n420), .b(n417), .O(n421));
  inv1   g348(.a(n420), .O(n422));
  nor2   g349(.a(n422), .b(n416), .O(n423));
  nor2   g350(.a(n423), .b(n421), .O(n424));
  nor2   g351(.a(n424), .b(n308), .O(n425));
  inv1   g352(.a(n424), .O(n426));
  nor2   g353(.a(n426), .b(n307), .O(n427));
  nor2   g354(.a(n427), .b(n425), .O(n428));
  inv1   g355(.a(n428), .O(n429));
  nor2   g356(.a(n429), .b(n414), .O(n430));
  nor2   g357(.a(n428), .b(n413), .O(n431));
  nor2   g358(.a(n431), .b(n430), .O(n432));
  inv1   g359(.a(n432), .O(n433));
  nor2   g360(.a(n433), .b(n406), .O(n434));
  inv1   g361(.a(n434), .O(n435));
  nor2   g362(.a(n435), .b(n380), .O(n436));
  inv1   g363(.a(n436), .O(n437));
  nor2   g364(.a(n437), .b(n277), .O(n438));
  inv1   g365(.a(n438), .O(n439));
  nor2   g366(.a(n439), .b(n137), .O(n440));
  nor2   g367(.a(n440), .b(n74), .O(n441));
  inv1   g368(.a(n440), .O(n442));
  nor2   g369(.a(n442), .b(G1gat), .O(n443));
  nor2   g370(.a(n443), .b(n441), .O(n444));
  inv1   g371(.a(n444), .O(G1324gat));
  nor2   g372(.a(n439), .b(n268), .O(n446));
  nor2   g373(.a(n446), .b(n248), .O(n447));
  inv1   g374(.a(n446), .O(n448));
  nor2   g375(.a(n448), .b(G8gat), .O(n449));
  nor2   g376(.a(n449), .b(n447), .O(n450));
  inv1   g377(.a(n450), .O(G1325gat));
  nor2   g378(.a(n439), .b(n232), .O(n452));
  nor2   g379(.a(n452), .b(n214), .O(n453));
  inv1   g380(.a(n452), .O(n454));
  nor2   g381(.a(n454), .b(G15gat), .O(n455));
  nor2   g382(.a(n455), .b(n453), .O(n456));
  inv1   g383(.a(n456), .O(G1326gat));
  nor2   g384(.a(n439), .b(n184), .O(n458));
  nor2   g385(.a(n458), .b(n167), .O(n459));
  inv1   g386(.a(n458), .O(n460));
  nor2   g387(.a(n460), .b(G22gat), .O(n461));
  nor2   g388(.a(n461), .b(n459), .O(n462));
  inv1   g389(.a(n462), .O(G1327gat));
  inv1   g390(.a(n406), .O(n464));
  nor2   g391(.a(n432), .b(n380), .O(n465));
  inv1   g392(.a(n465), .O(n466));
  nor2   g393(.a(n466), .b(n464), .O(n467));
  inv1   g394(.a(n467), .O(n468));
  nor2   g395(.a(n468), .b(n277), .O(n469));
  inv1   g396(.a(n469), .O(n470));
  nor2   g397(.a(n470), .b(n137), .O(n471));
  nor2   g398(.a(n471), .b(n119), .O(n472));
  inv1   g399(.a(n471), .O(n473));
  nor2   g400(.a(n473), .b(G29gat), .O(n474));
  nor2   g401(.a(n474), .b(n472), .O(n475));
  inv1   g402(.a(n475), .O(G1328gat));
  nor2   g403(.a(n470), .b(n268), .O(n477));
  nor2   g404(.a(n477), .b(n250), .O(n478));
  inv1   g405(.a(n477), .O(n479));
  nor2   g406(.a(n479), .b(G36gat), .O(n480));
  nor2   g407(.a(n480), .b(n478), .O(n481));
  inv1   g408(.a(n481), .O(G1329gat));
  nor2   g409(.a(n470), .b(n232), .O(n483));
  nor2   g410(.a(n483), .b(n216), .O(n484));
  inv1   g411(.a(n483), .O(n485));
  nor2   g412(.a(n485), .b(G43gat), .O(n486));
  nor2   g413(.a(n486), .b(n484), .O(n487));
  inv1   g414(.a(n487), .O(G1330gat));
  nor2   g415(.a(n470), .b(n184), .O(n489));
  nor2   g416(.a(n489), .b(n169), .O(n490));
  inv1   g417(.a(n489), .O(n491));
  nor2   g418(.a(n491), .b(G50gat), .O(n492));
  nor2   g419(.a(n492), .b(n490), .O(n493));
  inv1   g420(.a(n493), .O(G1331gat));
  inv1   g421(.a(n378), .O(n495));
  nor2   g422(.a(n495), .b(n327), .O(n496));
  inv1   g423(.a(n496), .O(n497));
  nor2   g424(.a(n497), .b(n435), .O(n498));
  inv1   g425(.a(n498), .O(n499));
  nor2   g426(.a(n499), .b(n277), .O(n500));
  inv1   g427(.a(n500), .O(n501));
  nor2   g428(.a(n501), .b(n137), .O(n502));
  nor2   g429(.a(n502), .b(n121), .O(n503));
  inv1   g430(.a(n502), .O(n504));
  nor2   g431(.a(n504), .b(G57gat), .O(n505));
  nor2   g432(.a(n505), .b(n503), .O(n506));
  inv1   g433(.a(n506), .O(G1332gat));
  nor2   g434(.a(n501), .b(n268), .O(n508));
  nor2   g435(.a(n508), .b(n242), .O(n509));
  inv1   g436(.a(n508), .O(n510));
  nor2   g437(.a(n510), .b(G64gat), .O(n511));
  nor2   g438(.a(n511), .b(n509), .O(n512));
  inv1   g439(.a(n512), .O(G1333gat));
  nor2   g440(.a(n501), .b(n232), .O(n514));
  nor2   g441(.a(n514), .b(n186), .O(n515));
  inv1   g442(.a(n514), .O(n516));
  nor2   g443(.a(n516), .b(G71gat), .O(n517));
  nor2   g444(.a(n517), .b(n515), .O(n518));
  inv1   g445(.a(n518), .O(G1334gat));
  nor2   g446(.a(n501), .b(n184), .O(n520));
  nor2   g447(.a(n520), .b(n139), .O(n521));
  inv1   g448(.a(n520), .O(n522));
  nor2   g449(.a(n522), .b(G78gat), .O(n523));
  nor2   g450(.a(n523), .b(n521), .O(n524));
  inv1   g451(.a(n524), .O(G1335gat));
  nor2   g452(.a(n497), .b(n432), .O(n526));
  inv1   g453(.a(n526), .O(n527));
  nor2   g454(.a(n527), .b(n464), .O(n528));
  inv1   g455(.a(n528), .O(n529));
  nor2   g456(.a(n529), .b(n277), .O(n530));
  inv1   g457(.a(n530), .O(n531));
  nor2   g458(.a(n531), .b(n137), .O(n532));
  nor2   g459(.a(n532), .b(n115), .O(n533));
  inv1   g460(.a(n532), .O(n534));
  nor2   g461(.a(n534), .b(G85gat), .O(n535));
  nor2   g462(.a(n535), .b(n533), .O(n536));
  inv1   g463(.a(n536), .O(G1336gat));
  nor2   g464(.a(n531), .b(n268), .O(n538));
  nor2   g465(.a(n538), .b(n244), .O(n539));
  inv1   g466(.a(n538), .O(n540));
  nor2   g467(.a(n540), .b(G92gat), .O(n541));
  nor2   g468(.a(n541), .b(n539), .O(n542));
  inv1   g469(.a(n542), .O(G1337gat));
  nor2   g470(.a(n531), .b(n232), .O(n544));
  nor2   g471(.a(n544), .b(n185), .O(n545));
  inv1   g472(.a(n544), .O(n546));
  nor2   g473(.a(n546), .b(G99gat), .O(n547));
  nor2   g474(.a(n547), .b(n545), .O(n548));
  inv1   g475(.a(n548), .O(G1338gat));
  nor2   g476(.a(n531), .b(n184), .O(n550));
  nor2   g477(.a(n550), .b(n138), .O(n551));
  inv1   g478(.a(n550), .O(n552));
  nor2   g479(.a(n552), .b(G106gat), .O(n553));
  nor2   g480(.a(n553), .b(n551), .O(n554));
  inv1   g481(.a(n554), .O(G1339gat));
  nor2   g482(.a(n432), .b(n464), .O(n556));
  nor2   g483(.a(n556), .b(n434), .O(n557));
  nor2   g484(.a(n378), .b(n327), .O(n558));
  inv1   g485(.a(n558), .O(n559));
  nor2   g486(.a(n559), .b(n557), .O(n560));
  nor2   g487(.a(n526), .b(n465), .O(n561));
  nor2   g488(.a(n561), .b(n406), .O(n562));
  nor2   g489(.a(n562), .b(n560), .O(n563));
  inv1   g490(.a(n233), .O(n564));
  nor2   g491(.a(n273), .b(n564), .O(n565));
  inv1   g492(.a(n565), .O(n566));
  nor2   g493(.a(n566), .b(n563), .O(n567));
  inv1   g494(.a(n567), .O(n568));
  nor2   g495(.a(n568), .b(n328), .O(n569));
  nor2   g496(.a(n569), .b(n75), .O(n570));
  inv1   g497(.a(n569), .O(n571));
  nor2   g498(.a(n571), .b(G113gat), .O(n572));
  nor2   g499(.a(n572), .b(n570), .O(n573));
  inv1   g500(.a(n573), .O(G1340gat));
  nor2   g501(.a(n568), .b(n495), .O(n575));
  nor2   g502(.a(n575), .b(n81), .O(n576));
  inv1   g503(.a(n575), .O(n577));
  nor2   g504(.a(n577), .b(G120gat), .O(n578));
  nor2   g505(.a(n578), .b(n576), .O(n579));
  inv1   g506(.a(n579), .O(G1341gat));
  nor2   g507(.a(n568), .b(n433), .O(n581));
  nor2   g508(.a(n581), .b(n83), .O(n582));
  inv1   g509(.a(n581), .O(n583));
  nor2   g510(.a(n583), .b(G127gat), .O(n584));
  nor2   g511(.a(n584), .b(n582), .O(n585));
  inv1   g512(.a(n585), .O(G1342gat));
  nor2   g513(.a(n568), .b(n464), .O(n587));
  nor2   g514(.a(n587), .b(n77), .O(n588));
  inv1   g515(.a(n587), .O(n589));
  nor2   g516(.a(n589), .b(G134gat), .O(n590));
  nor2   g517(.a(n590), .b(n588), .O(n591));
  inv1   g518(.a(n591), .O(G1343gat));
  inv1   g519(.a(n274), .O(n593));
  nor2   g520(.a(n593), .b(n184), .O(n594));
  inv1   g521(.a(n594), .O(n595));
  nor2   g522(.a(n595), .b(n563), .O(n596));
  inv1   g523(.a(n596), .O(n597));
  nor2   g524(.a(n597), .b(n328), .O(n598));
  nor2   g525(.a(n598), .b(n99), .O(n599));
  inv1   g526(.a(n598), .O(n600));
  nor2   g527(.a(n600), .b(G141gat), .O(n601));
  nor2   g528(.a(n601), .b(n599), .O(n602));
  inv1   g529(.a(n602), .O(G1344gat));
  nor2   g530(.a(n597), .b(n495), .O(n604));
  nor2   g531(.a(n604), .b(n105), .O(n605));
  inv1   g532(.a(n604), .O(n606));
  nor2   g533(.a(n606), .b(G148gat), .O(n607));
  nor2   g534(.a(n607), .b(n605), .O(n608));
  inv1   g535(.a(n608), .O(G1345gat));
  nor2   g536(.a(n597), .b(n433), .O(n610));
  nor2   g537(.a(n610), .b(n107), .O(n611));
  inv1   g538(.a(n610), .O(n612));
  nor2   g539(.a(n612), .b(G155gat), .O(n613));
  nor2   g540(.a(n613), .b(n611), .O(n614));
  inv1   g541(.a(n614), .O(G1346gat));
  nor2   g542(.a(n597), .b(n464), .O(n616));
  nor2   g543(.a(n616), .b(n101), .O(n617));
  inv1   g544(.a(n616), .O(n618));
  nor2   g545(.a(n618), .b(G162gat), .O(n619));
  nor2   g546(.a(n619), .b(n617), .O(n620));
  inv1   g547(.a(n620), .O(G1347gat));
  nor2   g548(.a(n270), .b(n564), .O(n622));
  inv1   g549(.a(n622), .O(n623));
  nor2   g550(.a(n623), .b(n563), .O(n624));
  inv1   g551(.a(n624), .O(n625));
  nor2   g552(.a(n625), .b(n328), .O(n626));
  nor2   g553(.a(n626), .b(n187), .O(n627));
  inv1   g554(.a(n626), .O(n628));
  nor2   g555(.a(n628), .b(G169gat), .O(n629));
  nor2   g556(.a(n629), .b(n627), .O(n630));
  inv1   g557(.a(n630), .O(G1348gat));
  nor2   g558(.a(n625), .b(n495), .O(n632));
  nor2   g559(.a(n632), .b(n193), .O(n633));
  inv1   g560(.a(n632), .O(n634));
  nor2   g561(.a(n634), .b(G176gat), .O(n635));
  nor2   g562(.a(n635), .b(n633), .O(n636));
  inv1   g563(.a(n636), .O(G1349gat));
  nor2   g564(.a(n625), .b(n433), .O(n638));
  nor2   g565(.a(n638), .b(n195), .O(n639));
  inv1   g566(.a(n638), .O(n640));
  nor2   g567(.a(n640), .b(G183gat), .O(n641));
  nor2   g568(.a(n641), .b(n639), .O(n642));
  inv1   g569(.a(n642), .O(G1350gat));
  nor2   g570(.a(n625), .b(n464), .O(n644));
  nor2   g571(.a(n644), .b(n189), .O(n645));
  inv1   g572(.a(n644), .O(n646));
  nor2   g573(.a(n646), .b(G190gat), .O(n647));
  nor2   g574(.a(n647), .b(n645), .O(n648));
  inv1   g575(.a(n648), .O(G1351gat));
  inv1   g576(.a(n271), .O(n650));
  nor2   g577(.a(n650), .b(n184), .O(n651));
  inv1   g578(.a(n651), .O(n652));
  nor2   g579(.a(n652), .b(n563), .O(n653));
  inv1   g580(.a(n653), .O(n654));
  nor2   g581(.a(n654), .b(n328), .O(n655));
  nor2   g582(.a(n655), .b(n140), .O(n656));
  inv1   g583(.a(n655), .O(n657));
  nor2   g584(.a(n657), .b(G197gat), .O(n658));
  nor2   g585(.a(n658), .b(n656), .O(n659));
  inv1   g586(.a(n659), .O(G1352gat));
  nor2   g587(.a(n654), .b(n495), .O(n661));
  nor2   g588(.a(n661), .b(n146), .O(n662));
  inv1   g589(.a(n661), .O(n663));
  nor2   g590(.a(n663), .b(G204gat), .O(n664));
  nor2   g591(.a(n664), .b(n662), .O(n665));
  inv1   g592(.a(n665), .O(G1353gat));
  nor2   g593(.a(n654), .b(n433), .O(n667));
  nor2   g594(.a(n667), .b(n148), .O(n668));
  inv1   g595(.a(n667), .O(n669));
  nor2   g596(.a(n669), .b(G211gat), .O(n670));
  nor2   g597(.a(n670), .b(n668), .O(n671));
  inv1   g598(.a(n671), .O(G1354gat));
  nor2   g599(.a(n654), .b(n464), .O(n673));
  nor2   g600(.a(n673), .b(n142), .O(n674));
  inv1   g601(.a(n673), .O(n675));
  nor2   g602(.a(n675), .b(G218gat), .O(n676));
  nor2   g603(.a(n676), .b(n674), .O(n677));
  inv1   g604(.a(n677), .O(G1355gat));
endmodule


