// Benchmark "c5315_blif" written by ABC on Sun Mar 24 18:39:14 2019

module c5315_blif  ( 
    G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37,
    G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79,
    G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106,
    G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140,
    G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173,
    G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209,
    G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251,
    G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293,
    G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338,
    G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389,
    G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523,
    G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691,
    G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717,
    G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115,
    G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612,
    G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921,
    G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636,
    G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626,
    G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623,
    G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000,
    G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802,
    G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826,
    G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742,
    G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843,
    G882, G767, G807, G658, G690  );
  input  G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34,
    G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76,
    G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103,
    G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121,
    G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137,
    G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170,
    G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206,
    G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248,
    G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292,
    G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335,
    G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386,
    G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514,
    G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690,
    G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552,
    G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115;
  output G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611,
    G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923,
    G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593,
    G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615,
    G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861,
    G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998,
    G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792,
    G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813,
    G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732,
    G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685,
    G688, G843, G882, G767, G807, G658, G690;
  wire n311, n312, n316, n317, n319, n321, n322, n324, n325, n326, n328,
    n329, n330, n332, n335, n336, n337, n338, n339, n340, n342, n343, n344,
    n345, n346, n348, n349, n351, n352, n353, n354, n355, n356, n357, n359,
    n360, n361, n362, n363, n364, n365, n367, n368, n369, n370, n371, n372,
    n373, n375, n376, n377, n378, n379, n380, n381, n383, n384, n385, n386,
    n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n487, n488, n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
    n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731, n732, n733, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n851, n852, n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
    n884, n885, n886, n888, n889, n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903, n904, n906, n907, n908, n909,
    n910, n911, n912, n913, n914, n915, n916, n917, n918, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n940, n941, n942, n943, n944, n945, n946, n947,
    n948, n949, n950, n951, n953, n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
    n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1028, n1029, n1030, n1031,
    n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1081, n1082, n1083, n1084,
    n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
    n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1153, n1154, n1155, n1156, n1157, n1158,
    n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
    n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
    n1189, n1190, n1191, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
    n1262, n1263, n1264, n1265, n1266, n1267, n1269, n1270, n1271, n1272,
    n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
    n1283, n1284, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
    n1349, n1350, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
    n1382, n1383, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
    n1393, n1394, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
    n1415, n1416, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
    n1448, n1449, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1485, n1486, n1487, n1489, n1490, n1491,
    n1492, n1493, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
    n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1523, n1524,
    n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1533, n1534, n1535,
    n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
    n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
    n1602, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
    n1613, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
    n1635, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
    n1657, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
    n1679, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
    n1712, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
    n1723, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
    n1745, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
    n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
    n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
    n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
    n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
    n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
    n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
    n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
    n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
    n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
    n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
    n1897, n1898, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
    n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
    n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
    n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
    n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
    n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
    n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
    n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
    n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
    n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
    n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
    n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
    n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
    n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
    n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
    n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2149,
    n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
    n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
    n2182;
  inv1   g0000(.a(G545), .O(G594));
  inv1   g0001(.a(G348), .O(G599));
  inv1   g0002(.a(G366), .O(G600));
  inv1   g0003(.a(G552), .O(G849));
  inv1   g0004(.a(G562), .O(G850));
  nor2   g0005(.a(G850), .b(G849), .O(G601));
  inv1   g0006(.a(G549), .O(G602));
  inv1   g0007(.a(G338), .O(G611));
  inv1   g0008(.a(G358), .O(G612));
  inv1   g0009(.a(G141), .O(n311));
  inv1   g0010(.a(G145), .O(n312));
  nor2   g0011(.a(n312), .b(n311), .O(G810));
  inv1   g0012(.a(G245), .O(G848));
  inv1   g0013(.a(G559), .O(G851));
  inv1   g0014(.a(G1), .O(n316));
  inv1   g0015(.a(G373), .O(n317));
  nor2   g0016(.a(n317), .b(n316), .O(G634));
  inv1   g0017(.a(G136), .O(n319));
  nor2   g0018(.a(G3173), .b(n319), .O(G815));
  inv1   g0019(.a(G27), .O(n321));
  nor2   g0020(.a(G2824), .b(n321), .O(n322));
  inv1   g0021(.a(n322), .O(G845));
  inv1   g0022(.a(G386), .O(n324));
  inv1   g0023(.a(G556), .O(n325));
  nor2   g0024(.a(n325), .b(n324), .O(n326));
  inv1   g0025(.a(n326), .O(G847));
  inv1   g0026(.a(G140), .O(n328));
  inv1   g0027(.a(G31), .O(n329));
  nor2   g0028(.a(n329), .b(n321), .O(n330));
  inv1   g0029(.a(n330), .O(G809));
  nor2   g0030(.a(G809), .b(n328), .O(n332));
  inv1   g0031(.a(n332), .O(G656));
  inv1   g0032(.a(G299), .O(G593));
  inv1   g0033(.a(G2358), .O(n335));
  nor2   g0034(.a(n335), .b(G87), .O(n336));
  nor2   g0035(.a(G2358), .b(G86), .O(n337));
  nor2   g0036(.a(n337), .b(G809), .O(n338));
  inv1   g0037(.a(n338), .O(n339));
  nor2   g0038(.a(n339), .b(n336), .O(n340));
  inv1   g0039(.a(n340), .O(G636));
  nor2   g0040(.a(n335), .b(G34), .O(n342));
  nor2   g0041(.a(G2358), .b(G88), .O(n343));
  nor2   g0042(.a(n343), .b(G809), .O(n344));
  inv1   g0043(.a(n344), .O(n345));
  nor2   g0044(.a(n345), .b(n342), .O(n346));
  inv1   g0045(.a(n346), .O(G704));
  inv1   g0046(.a(G83), .O(n348));
  nor2   g0047(.a(G809), .b(n348), .O(n349));
  inv1   g0048(.a(n349), .O(G820));
  inv1   g0049(.a(G25), .O(n351));
  nor2   g0050(.a(n335), .b(n351), .O(n352));
  inv1   g0051(.a(G24), .O(n353));
  nor2   g0052(.a(G2358), .b(n353), .O(n354));
  nor2   g0053(.a(n354), .b(G809), .O(n355));
  inv1   g0054(.a(n355), .O(n356));
  nor2   g0055(.a(n356), .b(n352), .O(n357));
  nor2   g0056(.a(n357), .b(n311), .O(G639));
  inv1   g0057(.a(G81), .O(n359));
  nor2   g0058(.a(n335), .b(n359), .O(n360));
  inv1   g0059(.a(G26), .O(n361));
  nor2   g0060(.a(G2358), .b(n361), .O(n362));
  nor2   g0061(.a(n362), .b(G809), .O(n363));
  inv1   g0062(.a(n363), .O(n364));
  nor2   g0063(.a(n364), .b(n360), .O(n365));
  nor2   g0064(.a(n365), .b(n311), .O(G673));
  inv1   g0065(.a(G23), .O(n367));
  nor2   g0066(.a(n335), .b(n367), .O(n368));
  inv1   g0067(.a(G79), .O(n369));
  nor2   g0068(.a(G2358), .b(n369), .O(n370));
  nor2   g0069(.a(n370), .b(G809), .O(n371));
  inv1   g0070(.a(n371), .O(n372));
  nor2   g0071(.a(n372), .b(n368), .O(n373));
  nor2   g0072(.a(n373), .b(n311), .O(G707));
  inv1   g0073(.a(G80), .O(n375));
  nor2   g0074(.a(n335), .b(n375), .O(n376));
  inv1   g0075(.a(G82), .O(n377));
  nor2   g0076(.a(G2358), .b(n377), .O(n378));
  nor2   g0077(.a(n378), .b(G809), .O(n379));
  inv1   g0078(.a(n379), .O(n380));
  nor2   g0079(.a(n380), .b(n376), .O(n381));
  nor2   g0080(.a(n381), .b(n311), .O(G715));
  inv1   g0081(.a(G341), .O(n383));
  inv1   g0082(.a(G3552), .O(n384));
  nor2   g0083(.a(n384), .b(n383), .O(n385));
  inv1   g0084(.a(G523), .O(n386));
  inv1   g0085(.a(G3550), .O(n387));
  nor2   g0086(.a(n387), .b(G341), .O(n388));
  nor2   g0087(.a(n388), .b(n386), .O(n389));
  inv1   g0088(.a(n389), .O(n390));
  nor2   g0089(.a(n390), .b(n385), .O(n391));
  nor2   g0090(.a(G3546), .b(n383), .O(n392));
  nor2   g0091(.a(G3548), .b(G341), .O(n393));
  nor2   g0092(.a(n393), .b(G523), .O(n394));
  inv1   g0093(.a(n394), .O(n395));
  nor2   g0094(.a(n395), .b(n392), .O(n396));
  nor2   g0095(.a(n396), .b(n391), .O(n397));
  inv1   g0096(.a(G351), .O(n398));
  nor2   g0097(.a(n384), .b(n398), .O(n399));
  inv1   g0098(.a(G534), .O(n400));
  nor2   g0099(.a(n387), .b(G351), .O(n401));
  nor2   g0100(.a(n401), .b(n400), .O(n402));
  inv1   g0101(.a(n402), .O(n403));
  nor2   g0102(.a(n403), .b(n399), .O(n404));
  nor2   g0103(.a(G3546), .b(n398), .O(n405));
  nor2   g0104(.a(G3548), .b(G351), .O(n406));
  nor2   g0105(.a(n406), .b(G534), .O(n407));
  inv1   g0106(.a(n407), .O(n408));
  nor2   g0107(.a(n408), .b(n405), .O(n409));
  nor2   g0108(.a(n409), .b(n404), .O(n410));
  inv1   g0109(.a(G324), .O(n411));
  nor2   g0110(.a(n384), .b(n411), .O(n412));
  inv1   g0111(.a(G503), .O(n413));
  nor2   g0112(.a(n387), .b(G324), .O(n414));
  nor2   g0113(.a(n414), .b(n413), .O(n415));
  inv1   g0114(.a(n415), .O(n416));
  nor2   g0115(.a(n416), .b(n412), .O(n417));
  nor2   g0116(.a(G3546), .b(n411), .O(n418));
  nor2   g0117(.a(G3548), .b(G324), .O(n419));
  nor2   g0118(.a(n419), .b(G503), .O(n420));
  inv1   g0119(.a(n420), .O(n421));
  nor2   g0120(.a(n421), .b(n418), .O(n422));
  nor2   g0121(.a(n422), .b(n417), .O(n423));
  nor2   g0122(.a(n423), .b(n410), .O(n424));
  inv1   g0123(.a(n424), .O(n425));
  nor2   g0124(.a(n425), .b(n397), .O(n426));
  inv1   g0125(.a(n426), .O(n427));
  inv1   g0126(.a(G248), .O(n428));
  inv1   g0127(.a(G302), .O(n429));
  nor2   g0128(.a(n429), .b(n428), .O(n430));
  inv1   g0129(.a(G251), .O(n431));
  nor2   g0130(.a(G302), .b(n431), .O(n432));
  nor2   g0131(.a(n432), .b(n430), .O(n433));
  inv1   g0132(.a(G308), .O(n434));
  nor2   g0133(.a(n434), .b(G248), .O(n435));
  inv1   g0134(.a(G479), .O(n436));
  nor2   g0135(.a(G308), .b(G251), .O(n437));
  nor2   g0136(.a(n437), .b(n436), .O(n438));
  inv1   g0137(.a(n438), .O(n439));
  nor2   g0138(.a(n439), .b(n435), .O(n440));
  inv1   g0139(.a(G242), .O(n441));
  nor2   g0140(.a(n434), .b(n441), .O(n442));
  inv1   g0141(.a(G254), .O(n443));
  nor2   g0142(.a(G308), .b(n443), .O(n444));
  nor2   g0143(.a(n444), .b(G479), .O(n445));
  inv1   g0144(.a(n445), .O(n446));
  nor2   g0145(.a(n446), .b(n442), .O(n447));
  nor2   g0146(.a(n447), .b(n440), .O(n448));
  nor2   g0147(.a(n448), .b(n433), .O(n449));
  inv1   g0148(.a(n449), .O(n450));
  inv1   g0149(.a(G316), .O(n451));
  nor2   g0150(.a(n451), .b(G248), .O(n452));
  inv1   g0151(.a(G490), .O(n453));
  nor2   g0152(.a(G316), .b(G251), .O(n454));
  nor2   g0153(.a(n454), .b(n453), .O(n455));
  inv1   g0154(.a(n455), .O(n456));
  nor2   g0155(.a(n456), .b(n452), .O(n457));
  nor2   g0156(.a(n451), .b(n441), .O(n458));
  nor2   g0157(.a(G316), .b(n443), .O(n459));
  nor2   g0158(.a(n459), .b(G490), .O(n460));
  inv1   g0159(.a(n460), .O(n461));
  nor2   g0160(.a(n461), .b(n458), .O(n462));
  nor2   g0161(.a(n462), .b(n457), .O(n463));
  inv1   g0162(.a(G361), .O(n464));
  nor2   g0163(.a(n464), .b(n428), .O(n465));
  nor2   g0164(.a(G361), .b(n431), .O(n466));
  nor2   g0165(.a(n466), .b(n465), .O(n467));
  inv1   g0166(.a(G293), .O(n468));
  nor2   g0167(.a(n468), .b(n441), .O(n469));
  nor2   g0168(.a(G293), .b(n443), .O(n470));
  nor2   g0169(.a(n470), .b(n469), .O(n471));
  inv1   g0170(.a(n471), .O(n472));
  nor2   g0171(.a(n472), .b(n467), .O(n473));
  inv1   g0172(.a(n473), .O(n474));
  inv1   g0173(.a(G514), .O(n475));
  nor2   g0174(.a(G3552), .b(n475), .O(n476));
  inv1   g0175(.a(G3546), .O(n477));
  nor2   g0176(.a(n477), .b(G514), .O(n478));
  nor2   g0177(.a(n478), .b(n476), .O(n479));
  nor2   g0178(.a(n479), .b(n474), .O(n480));
  inv1   g0179(.a(n480), .O(n481));
  nor2   g0180(.a(n481), .b(n463), .O(n482));
  inv1   g0181(.a(n482), .O(n483));
  nor2   g0182(.a(n483), .b(n450), .O(n484));
  inv1   g0183(.a(n484), .O(n485));
  nor2   g0184(.a(n485), .b(n427), .O(G598));
  inv1   g0185(.a(G265), .O(n487));
  nor2   g0186(.a(n384), .b(n487), .O(n488));
  inv1   g0187(.a(G400), .O(n489));
  nor2   g0188(.a(n387), .b(G265), .O(n490));
  nor2   g0189(.a(n490), .b(n489), .O(n491));
  inv1   g0190(.a(n491), .O(n492));
  nor2   g0191(.a(n492), .b(n488), .O(n493));
  nor2   g0192(.a(G3546), .b(n487), .O(n494));
  nor2   g0193(.a(G3548), .b(G265), .O(n495));
  nor2   g0194(.a(n495), .b(G400), .O(n496));
  inv1   g0195(.a(n496), .O(n497));
  nor2   g0196(.a(n497), .b(n494), .O(n498));
  nor2   g0197(.a(n498), .b(n493), .O(n499));
  inv1   g0198(.a(G210), .O(n500));
  nor2   g0199(.a(G3546), .b(n500), .O(n501));
  nor2   g0200(.a(G3548), .b(G210), .O(n502));
  nor2   g0201(.a(n502), .b(G457), .O(n503));
  inv1   g0202(.a(n503), .O(n504));
  nor2   g0203(.a(n504), .b(n501), .O(n505));
  inv1   g0204(.a(G457), .O(n506));
  nor2   g0205(.a(n506), .b(n500), .O(n507));
  inv1   g0206(.a(n507), .O(n508));
  nor2   g0207(.a(n508), .b(G3552), .O(n509));
  nor2   g0208(.a(n506), .b(G210), .O(n510));
  inv1   g0209(.a(n510), .O(n511));
  nor2   g0210(.a(n511), .b(G3550), .O(n512));
  nor2   g0211(.a(n512), .b(n509), .O(n513));
  inv1   g0212(.a(n513), .O(n514));
  nor2   g0213(.a(n514), .b(n505), .O(n515));
  inv1   g0214(.a(G273), .O(n516));
  nor2   g0215(.a(n384), .b(n516), .O(n517));
  inv1   g0216(.a(G411), .O(n518));
  nor2   g0217(.a(n387), .b(G273), .O(n519));
  nor2   g0218(.a(n519), .b(n518), .O(n520));
  inv1   g0219(.a(n520), .O(n521));
  nor2   g0220(.a(n521), .b(n517), .O(n522));
  nor2   g0221(.a(G3546), .b(n516), .O(n523));
  nor2   g0222(.a(G3548), .b(G273), .O(n524));
  nor2   g0223(.a(n524), .b(G411), .O(n525));
  inv1   g0224(.a(n525), .O(n526));
  nor2   g0225(.a(n526), .b(n523), .O(n527));
  nor2   g0226(.a(n527), .b(n522), .O(n528));
  nor2   g0227(.a(n528), .b(n515), .O(n529));
  inv1   g0228(.a(n529), .O(n530));
  nor2   g0229(.a(n530), .b(n499), .O(n531));
  inv1   g0230(.a(n531), .O(n532));
  inv1   g0231(.a(G226), .O(n533));
  nor2   g0232(.a(G3546), .b(n533), .O(n534));
  nor2   g0233(.a(G3548), .b(G226), .O(n535));
  nor2   g0234(.a(n535), .b(G422), .O(n536));
  inv1   g0235(.a(n536), .O(n537));
  nor2   g0236(.a(n537), .b(n534), .O(n538));
  inv1   g0237(.a(G422), .O(n539));
  nor2   g0238(.a(n539), .b(n533), .O(n540));
  inv1   g0239(.a(n540), .O(n541));
  nor2   g0240(.a(n541), .b(G3552), .O(n542));
  nor2   g0241(.a(n539), .b(G226), .O(n543));
  inv1   g0242(.a(n543), .O(n544));
  nor2   g0243(.a(n544), .b(G3550), .O(n545));
  nor2   g0244(.a(n545), .b(n542), .O(n546));
  inv1   g0245(.a(n546), .O(n547));
  nor2   g0246(.a(n547), .b(n538), .O(n548));
  inv1   g0247(.a(G281), .O(n549));
  nor2   g0248(.a(n384), .b(n549), .O(n550));
  inv1   g0249(.a(G374), .O(n551));
  nor2   g0250(.a(n387), .b(G281), .O(n552));
  nor2   g0251(.a(n552), .b(n551), .O(n553));
  inv1   g0252(.a(n553), .O(n554));
  nor2   g0253(.a(n554), .b(n550), .O(n555));
  nor2   g0254(.a(G3546), .b(n549), .O(n556));
  nor2   g0255(.a(G3548), .b(G281), .O(n557));
  nor2   g0256(.a(n557), .b(G374), .O(n558));
  inv1   g0257(.a(n558), .O(n559));
  nor2   g0258(.a(n559), .b(n556), .O(n560));
  nor2   g0259(.a(n560), .b(n555), .O(n561));
  nor2   g0260(.a(n561), .b(n548), .O(n562));
  inv1   g0261(.a(n562), .O(n563));
  inv1   g0262(.a(G257), .O(n564));
  nor2   g0263(.a(n384), .b(n564), .O(n565));
  inv1   g0264(.a(G389), .O(n566));
  nor2   g0265(.a(n387), .b(G257), .O(n567));
  nor2   g0266(.a(n567), .b(n566), .O(n568));
  inv1   g0267(.a(n568), .O(n569));
  nor2   g0268(.a(n569), .b(n565), .O(n570));
  nor2   g0269(.a(G3546), .b(n564), .O(n571));
  nor2   g0270(.a(G3548), .b(G257), .O(n572));
  nor2   g0271(.a(n572), .b(G389), .O(n573));
  inv1   g0272(.a(n573), .O(n574));
  nor2   g0273(.a(n574), .b(n571), .O(n575));
  nor2   g0274(.a(n575), .b(n570), .O(n576));
  inv1   g0275(.a(G234), .O(n577));
  nor2   g0276(.a(G3546), .b(n577), .O(n578));
  nor2   g0277(.a(G3548), .b(G234), .O(n579));
  nor2   g0278(.a(n579), .b(G435), .O(n580));
  inv1   g0279(.a(n580), .O(n581));
  nor2   g0280(.a(n581), .b(n578), .O(n582));
  inv1   g0281(.a(G435), .O(n583));
  nor2   g0282(.a(n583), .b(n577), .O(n584));
  inv1   g0283(.a(n584), .O(n585));
  nor2   g0284(.a(n585), .b(G3552), .O(n586));
  nor2   g0285(.a(n583), .b(G234), .O(n587));
  inv1   g0286(.a(n587), .O(n588));
  nor2   g0287(.a(n588), .b(G3550), .O(n589));
  nor2   g0288(.a(n589), .b(n586), .O(n590));
  inv1   g0289(.a(n590), .O(n591));
  nor2   g0290(.a(n591), .b(n582), .O(n592));
  nor2   g0291(.a(n592), .b(n576), .O(n593));
  inv1   g0292(.a(n593), .O(n594));
  inv1   g0293(.a(G206), .O(n595));
  nor2   g0294(.a(G248), .b(n595), .O(n596));
  inv1   g0295(.a(G446), .O(n597));
  nor2   g0296(.a(G251), .b(G206), .O(n598));
  nor2   g0297(.a(n598), .b(n597), .O(n599));
  inv1   g0298(.a(n599), .O(n600));
  nor2   g0299(.a(n600), .b(n596), .O(n601));
  nor2   g0300(.a(n441), .b(n595), .O(n602));
  nor2   g0301(.a(n443), .b(G206), .O(n603));
  nor2   g0302(.a(n603), .b(G446), .O(n604));
  inv1   g0303(.a(n604), .O(n605));
  nor2   g0304(.a(n605), .b(n602), .O(n606));
  nor2   g0305(.a(n606), .b(n601), .O(n607));
  inv1   g0306(.a(G218), .O(n608));
  nor2   g0307(.a(G3546), .b(n608), .O(n609));
  nor2   g0308(.a(G3548), .b(G218), .O(n610));
  nor2   g0309(.a(n610), .b(G468), .O(n611));
  inv1   g0310(.a(n611), .O(n612));
  nor2   g0311(.a(n612), .b(n609), .O(n613));
  inv1   g0312(.a(G468), .O(n614));
  nor2   g0313(.a(n614), .b(n608), .O(n615));
  inv1   g0314(.a(n615), .O(n616));
  nor2   g0315(.a(n616), .b(G3552), .O(n617));
  nor2   g0316(.a(n614), .b(G218), .O(n618));
  inv1   g0317(.a(n618), .O(n619));
  nor2   g0318(.a(n619), .b(G3550), .O(n620));
  nor2   g0319(.a(n620), .b(n617), .O(n621));
  inv1   g0320(.a(n621), .O(n622));
  nor2   g0321(.a(n622), .b(n613), .O(n623));
  nor2   g0322(.a(n623), .b(n607), .O(n624));
  inv1   g0323(.a(n624), .O(n625));
  nor2   g0324(.a(n625), .b(n594), .O(n626));
  inv1   g0325(.a(n626), .O(n627));
  nor2   g0326(.a(n627), .b(n563), .O(n628));
  inv1   g0327(.a(n628), .O(n629));
  nor2   g0328(.a(n629), .b(n532), .O(G610));
  nor2   g0329(.a(G335), .b(n577), .O(n631));
  inv1   g0330(.a(G241), .O(n632));
  inv1   g0331(.a(G335), .O(n633));
  nor2   g0332(.a(n633), .b(n632), .O(n634));
  nor2   g0333(.a(n634), .b(n631), .O(n635));
  nor2   g0334(.a(n635), .b(n583), .O(n636));
  inv1   g0335(.a(n635), .O(n637));
  nor2   g0336(.a(n637), .b(G435), .O(n638));
  nor2   g0337(.a(n638), .b(n636), .O(n639));
  inv1   g0338(.a(n639), .O(n640));
  nor2   g0339(.a(G335), .b(n516), .O(n641));
  inv1   g0340(.a(G280), .O(n642));
  nor2   g0341(.a(n633), .b(n642), .O(n643));
  nor2   g0342(.a(n643), .b(n641), .O(n644));
  nor2   g0343(.a(n644), .b(n518), .O(n645));
  inv1   g0344(.a(n644), .O(n646));
  nor2   g0345(.a(n646), .b(G411), .O(n647));
  nor2   g0346(.a(n647), .b(n645), .O(n648));
  inv1   g0347(.a(n648), .O(n649));
  nor2   g0348(.a(G335), .b(n487), .O(n650));
  inv1   g0349(.a(G272), .O(n651));
  nor2   g0350(.a(n633), .b(n651), .O(n652));
  nor2   g0351(.a(n652), .b(n650), .O(n653));
  nor2   g0352(.a(n653), .b(n489), .O(n654));
  inv1   g0353(.a(n653), .O(n655));
  nor2   g0354(.a(n655), .b(G400), .O(n656));
  nor2   g0355(.a(n656), .b(n654), .O(n657));
  inv1   g0356(.a(n657), .O(n658));
  nor2   g0357(.a(n658), .b(n649), .O(n659));
  inv1   g0358(.a(n659), .O(n660));
  nor2   g0359(.a(G335), .b(n549), .O(n661));
  inv1   g0360(.a(G288), .O(n662));
  nor2   g0361(.a(n633), .b(n662), .O(n663));
  nor2   g0362(.a(n663), .b(n661), .O(n664));
  inv1   g0363(.a(n664), .O(n665));
  nor2   g0364(.a(n665), .b(G374), .O(n666));
  nor2   g0365(.a(n666), .b(n660), .O(n667));
  inv1   g0366(.a(n667), .O(n668));
  nor2   g0367(.a(n664), .b(n551), .O(n669));
  nor2   g0368(.a(G335), .b(n564), .O(n670));
  inv1   g0369(.a(G264), .O(n671));
  nor2   g0370(.a(n633), .b(n671), .O(n672));
  nor2   g0371(.a(n672), .b(n670), .O(n673));
  nor2   g0372(.a(n673), .b(n566), .O(n674));
  inv1   g0373(.a(n673), .O(n675));
  nor2   g0374(.a(n675), .b(G389), .O(n676));
  nor2   g0375(.a(n676), .b(n674), .O(n677));
  inv1   g0376(.a(n677), .O(n678));
  nor2   g0377(.a(n678), .b(n669), .O(n679));
  inv1   g0378(.a(n679), .O(n680));
  nor2   g0379(.a(n680), .b(n668), .O(n681));
  inv1   g0380(.a(n681), .O(n682));
  nor2   g0381(.a(n682), .b(n640), .O(n683));
  inv1   g0382(.a(n683), .O(n684));
  nor2   g0383(.a(G335), .b(n500), .O(n685));
  inv1   g0384(.a(G217), .O(n686));
  nor2   g0385(.a(n633), .b(n686), .O(n687));
  nor2   g0386(.a(n687), .b(n685), .O(n688));
  nor2   g0387(.a(n688), .b(n506), .O(n689));
  inv1   g0388(.a(n688), .O(n690));
  nor2   g0389(.a(n690), .b(G457), .O(n691));
  nor2   g0390(.a(n691), .b(n689), .O(n692));
  inv1   g0391(.a(n692), .O(n693));
  nor2   g0392(.a(G335), .b(n533), .O(n694));
  inv1   g0393(.a(G233), .O(n695));
  nor2   g0394(.a(n633), .b(n695), .O(n696));
  nor2   g0395(.a(n696), .b(n694), .O(n697));
  inv1   g0396(.a(n697), .O(n698));
  nor2   g0397(.a(n698), .b(G422), .O(n699));
  nor2   g0398(.a(G335), .b(n608), .O(n700));
  inv1   g0399(.a(G225), .O(n701));
  nor2   g0400(.a(n633), .b(n701), .O(n702));
  nor2   g0401(.a(n702), .b(n700), .O(n703));
  nor2   g0402(.a(n703), .b(n614), .O(n704));
  inv1   g0403(.a(n703), .O(n705));
  nor2   g0404(.a(n705), .b(G468), .O(n706));
  nor2   g0405(.a(n706), .b(n704), .O(n707));
  inv1   g0406(.a(n707), .O(n708));
  nor2   g0407(.a(n708), .b(n699), .O(n709));
  inv1   g0408(.a(n699), .O(n710));
  nor2   g0409(.a(n707), .b(n710), .O(n711));
  nor2   g0410(.a(n711), .b(n709), .O(n712));
  nor2   g0411(.a(n712), .b(n693), .O(n713));
  inv1   g0412(.a(n713), .O(n714));
  nor2   g0413(.a(G335), .b(n595), .O(n715));
  inv1   g0414(.a(G209), .O(n716));
  nor2   g0415(.a(n633), .b(n716), .O(n717));
  nor2   g0416(.a(n717), .b(n715), .O(n718));
  nor2   g0417(.a(n718), .b(n597), .O(n719));
  inv1   g0418(.a(n718), .O(n720));
  nor2   g0419(.a(n720), .b(G446), .O(n721));
  nor2   g0420(.a(n721), .b(n719), .O(n722));
  inv1   g0421(.a(n722), .O(n723));
  nor2   g0422(.a(n697), .b(n539), .O(n724));
  inv1   g0423(.a(n724), .O(n725));
  nor2   g0424(.a(n725), .b(n708), .O(n726));
  nor2   g0425(.a(n724), .b(n707), .O(n727));
  nor2   g0426(.a(n727), .b(n726), .O(n728));
  inv1   g0427(.a(n728), .O(n729));
  nor2   g0428(.a(n729), .b(n723), .O(n730));
  inv1   g0429(.a(n730), .O(n731));
  nor2   g0430(.a(n731), .b(n714), .O(n732));
  inv1   g0431(.a(n732), .O(n733));
  nor2   g0432(.a(n733), .b(n684), .O(G588));
  nor2   g0433(.a(G332), .b(n429), .O(n735));
  inv1   g0434(.a(G307), .O(n736));
  inv1   g0435(.a(G332), .O(n737));
  nor2   g0436(.a(n737), .b(n736), .O(n738));
  nor2   g0437(.a(n738), .b(n735), .O(n739));
  inv1   g0438(.a(n739), .O(n740));
  nor2   g0439(.a(G332), .b(n468), .O(n741));
  nor2   g0440(.a(n737), .b(G593), .O(n742));
  nor2   g0441(.a(n742), .b(n741), .O(n743));
  inv1   g0442(.a(n743), .O(n744));
  nor2   g0443(.a(n744), .b(n740), .O(n745));
  inv1   g0444(.a(n745), .O(n746));
  nor2   g0445(.a(G332), .b(n451), .O(n747));
  inv1   g0446(.a(G323), .O(n748));
  nor2   g0447(.a(n737), .b(n748), .O(n749));
  nor2   g0448(.a(n749), .b(n747), .O(n750));
  nor2   g0449(.a(n750), .b(n453), .O(n751));
  inv1   g0450(.a(n750), .O(n752));
  nor2   g0451(.a(n752), .b(G490), .O(n753));
  nor2   g0452(.a(n753), .b(n751), .O(n754));
  inv1   g0453(.a(n754), .O(n755));
  nor2   g0454(.a(G332), .b(n434), .O(n756));
  inv1   g0455(.a(G315), .O(n757));
  nor2   g0456(.a(n737), .b(n757), .O(n758));
  nor2   g0457(.a(n758), .b(n756), .O(n759));
  nor2   g0458(.a(n759), .b(n436), .O(n760));
  inv1   g0459(.a(n759), .O(n761));
  nor2   g0460(.a(n761), .b(G479), .O(n762));
  nor2   g0461(.a(n762), .b(n760), .O(n763));
  inv1   g0462(.a(n763), .O(n764));
  nor2   g0463(.a(n764), .b(n755), .O(n765));
  inv1   g0464(.a(n765), .O(n766));
  nor2   g0465(.a(n766), .b(n746), .O(n767));
  inv1   g0466(.a(n767), .O(n768));
  nor2   g0467(.a(n383), .b(G332), .O(n769));
  nor2   g0468(.a(G599), .b(n737), .O(n770));
  nor2   g0469(.a(n770), .b(n769), .O(n771));
  nor2   g0470(.a(n771), .b(n386), .O(n772));
  inv1   g0471(.a(n771), .O(n773));
  nor2   g0472(.a(n773), .b(G523), .O(n774));
  nor2   g0473(.a(n774), .b(n772), .O(n775));
  inv1   g0474(.a(n775), .O(n776));
  nor2   g0475(.a(n398), .b(G332), .O(n777));
  nor2   g0476(.a(G612), .b(n737), .O(n778));
  nor2   g0477(.a(n778), .b(n777), .O(n779));
  inv1   g0478(.a(n779), .O(n780));
  nor2   g0479(.a(n780), .b(G534), .O(n781));
  nor2   g0480(.a(n779), .b(n400), .O(n782));
  nor2   g0481(.a(n782), .b(n781), .O(n783));
  inv1   g0482(.a(n783), .O(n784));
  nor2   g0483(.a(n464), .b(G332), .O(n785));
  nor2   g0484(.a(G600), .b(n737), .O(n786));
  nor2   g0485(.a(n786), .b(n785), .O(n787));
  inv1   g0486(.a(n787), .O(n788));
  nor2   g0487(.a(n788), .b(n784), .O(n789));
  inv1   g0488(.a(n789), .O(n790));
  nor2   g0489(.a(n790), .b(n776), .O(n791));
  inv1   g0490(.a(n791), .O(n792));
  nor2   g0491(.a(G338), .b(n737), .O(n793));
  inv1   g0492(.a(n793), .O(n794));
  nor2   g0493(.a(n794), .b(G514), .O(n795));
  nor2   g0494(.a(n795), .b(n792), .O(n796));
  inv1   g0495(.a(n796), .O(n797));
  nor2   g0496(.a(n737), .b(G331), .O(n798));
  nor2   g0497(.a(G332), .b(G324), .O(n799));
  nor2   g0498(.a(n799), .b(n798), .O(n800));
  inv1   g0499(.a(n800), .O(n801));
  nor2   g0500(.a(n801), .b(n413), .O(n802));
  nor2   g0501(.a(n800), .b(G503), .O(n803));
  nor2   g0502(.a(n803), .b(n802), .O(n804));
  inv1   g0503(.a(n804), .O(n805));
  nor2   g0504(.a(n793), .b(n475), .O(n806));
  nor2   g0505(.a(n789), .b(n781), .O(n807));
  nor2   g0506(.a(n807), .b(n772), .O(n808));
  nor2   g0507(.a(n808), .b(n774), .O(n809));
  nor2   g0508(.a(n809), .b(n806), .O(n810));
  inv1   g0509(.a(n809), .O(n811));
  nor2   g0510(.a(n811), .b(n795), .O(n812));
  nor2   g0511(.a(n812), .b(n810), .O(n813));
  nor2   g0512(.a(n813), .b(n805), .O(n814));
  inv1   g0513(.a(n814), .O(n815));
  nor2   g0514(.a(n815), .b(n797), .O(n816));
  inv1   g0515(.a(n816), .O(n817));
  nor2   g0516(.a(n817), .b(n768), .O(G615));
  nor2   g0517(.a(G316), .b(n434), .O(n819));
  nor2   g0518(.a(n451), .b(G308), .O(n820));
  nor2   g0519(.a(n820), .b(n819), .O(n821));
  inv1   g0520(.a(n821), .O(n822));
  nor2   g0521(.a(G351), .b(n383), .O(n823));
  nor2   g0522(.a(n398), .b(G341), .O(n824));
  nor2   g0523(.a(n824), .b(n823), .O(n825));
  inv1   g0524(.a(n825), .O(n826));
  nor2   g0525(.a(n826), .b(n468), .O(n827));
  nor2   g0526(.a(n825), .b(G293), .O(n828));
  nor2   g0527(.a(n828), .b(n827), .O(n829));
  inv1   g0528(.a(n829), .O(n830));
  nor2   g0529(.a(G369), .b(n464), .O(n831));
  inv1   g0530(.a(G369), .O(n832));
  nor2   g0531(.a(n832), .b(G361), .O(n833));
  nor2   g0532(.a(n833), .b(n831), .O(n834));
  inv1   g0533(.a(n834), .O(n835));
  nor2   g0534(.a(G324), .b(n429), .O(n836));
  nor2   g0535(.a(n411), .b(G302), .O(n837));
  nor2   g0536(.a(n837), .b(n836), .O(n838));
  inv1   g0537(.a(n838), .O(n839));
  nor2   g0538(.a(n839), .b(n835), .O(n840));
  nor2   g0539(.a(n838), .b(n834), .O(n841));
  nor2   g0540(.a(n841), .b(n840), .O(n842));
  nor2   g0541(.a(n842), .b(n830), .O(n843));
  inv1   g0542(.a(n842), .O(n844));
  nor2   g0543(.a(n844), .b(n829), .O(n845));
  nor2   g0544(.a(n845), .b(n843), .O(n846));
  inv1   g0545(.a(n846), .O(n847));
  nor2   g0546(.a(n847), .b(n822), .O(n848));
  nor2   g0547(.a(n846), .b(n821), .O(n849));
  nor2   g0548(.a(n849), .b(n848), .O(G1002));
  nor2   g0549(.a(G257), .b(n577), .O(n851));
  nor2   g0550(.a(n564), .b(G234), .O(n852));
  nor2   g0551(.a(n852), .b(n851), .O(n853));
  inv1   g0552(.a(n853), .O(n854));
  nor2   g0553(.a(G273), .b(n487), .O(n855));
  nor2   g0554(.a(n516), .b(G265), .O(n856));
  nor2   g0555(.a(n856), .b(n855), .O(n857));
  inv1   g0556(.a(n857), .O(n858));
  nor2   g0557(.a(n858), .b(n595), .O(n859));
  nor2   g0558(.a(n857), .b(G206), .O(n860));
  nor2   g0559(.a(n860), .b(n859), .O(n861));
  nor2   g0560(.a(n861), .b(n854), .O(n862));
  inv1   g0561(.a(n861), .O(n863));
  nor2   g0562(.a(n863), .b(n853), .O(n864));
  nor2   g0563(.a(n864), .b(n862), .O(n865));
  inv1   g0564(.a(n865), .O(n866));
  inv1   g0565(.a(G289), .O(n867));
  nor2   g0566(.a(G281), .b(G210), .O(n868));
  nor2   g0567(.a(n549), .b(n500), .O(n869));
  nor2   g0568(.a(n869), .b(n868), .O(n870));
  inv1   g0569(.a(n870), .O(n871));
  nor2   g0570(.a(n871), .b(n867), .O(n872));
  nor2   g0571(.a(n870), .b(G289), .O(n873));
  nor2   g0572(.a(n873), .b(n872), .O(n874));
  inv1   g0573(.a(n874), .O(n875));
  nor2   g0574(.a(G226), .b(n608), .O(n876));
  nor2   g0575(.a(n533), .b(G218), .O(n877));
  nor2   g0576(.a(n877), .b(n876), .O(n878));
  nor2   g0577(.a(n878), .b(n875), .O(n879));
  inv1   g0578(.a(n878), .O(n880));
  nor2   g0579(.a(n880), .b(n874), .O(n881));
  nor2   g0580(.a(n881), .b(n879), .O(n882));
  inv1   g0581(.a(n882), .O(n883));
  nor2   g0582(.a(n883), .b(n866), .O(n884));
  nor2   g0583(.a(n882), .b(n865), .O(n885));
  nor2   g0584(.a(n885), .b(n884), .O(n886));
  inv1   g0585(.a(n886), .O(G1004));
  inv1   g0586(.a(n669), .O(n888));
  nor2   g0587(.a(n888), .b(n660), .O(n889));
  nor2   g0588(.a(n654), .b(n645), .O(n890));
  nor2   g0589(.a(n890), .b(n656), .O(n891));
  nor2   g0590(.a(n891), .b(n889), .O(n892));
  nor2   g0591(.a(n892), .b(n676), .O(n893));
  nor2   g0592(.a(n893), .b(n674), .O(n894));
  nor2   g0593(.a(n894), .b(n638), .O(n895));
  nor2   g0594(.a(n895), .b(n636), .O(n896));
  nor2   g0595(.a(n896), .b(n733), .O(n897));
  nor2   g0596(.a(n726), .b(n704), .O(n898));
  nor2   g0597(.a(n898), .b(n691), .O(n899));
  nor2   g0598(.a(n899), .b(n689), .O(n900));
  nor2   g0599(.a(n900), .b(n721), .O(n901));
  nor2   g0600(.a(n901), .b(n719), .O(n902));
  inv1   g0601(.a(n902), .O(n903));
  nor2   g0602(.a(n903), .b(n897), .O(n904));
  inv1   g0603(.a(n904), .O(G591));
  nor2   g0604(.a(n806), .b(n802), .O(n906));
  inv1   g0605(.a(n906), .O(n907));
  nor2   g0606(.a(n907), .b(n812), .O(n908));
  nor2   g0607(.a(n908), .b(n803), .O(n909));
  inv1   g0608(.a(n909), .O(n910));
  nor2   g0609(.a(n910), .b(n768), .O(n911));
  inv1   g0610(.a(n751), .O(n912));
  nor2   g0611(.a(n764), .b(n912), .O(n913));
  nor2   g0612(.a(n913), .b(n760), .O(n914));
  inv1   g0613(.a(n914), .O(n915));
  nor2   g0614(.a(n915), .b(n746), .O(n916));
  inv1   g0615(.a(n916), .O(n917));
  nor2   g0616(.a(n917), .b(n911), .O(n918));
  inv1   g0617(.a(n918), .O(G618));
  nor2   g0618(.a(n788), .b(G54), .O(n920));
  inv1   g0619(.a(G54), .O(n921));
  nor2   g0620(.a(n787), .b(n921), .O(n922));
  nor2   g0621(.a(n922), .b(n920), .O(n923));
  inv1   g0622(.a(G4091), .O(n924));
  nor2   g0623(.a(G4092), .b(n924), .O(n925));
  inv1   g0624(.a(n925), .O(n926));
  nor2   g0625(.a(n926), .b(n923), .O(n927));
  inv1   g0626(.a(n467), .O(n928));
  nor2   g0627(.a(G4092), .b(G4091), .O(n929));
  inv1   g0628(.a(n929), .O(n930));
  nor2   g0629(.a(n930), .b(n928), .O(n931));
  inv1   g0630(.a(G131), .O(n932));
  inv1   g0631(.a(G4092), .O(n933));
  nor2   g0632(.a(n933), .b(G4091), .O(n934));
  inv1   g0633(.a(n934), .O(n935));
  nor2   g0634(.a(n935), .b(n932), .O(n936));
  nor2   g0635(.a(n936), .b(n931), .O(n937));
  inv1   g0636(.a(n937), .O(n938));
  nor2   g0637(.a(n938), .b(n927), .O(G822));
  nor2   g0638(.a(n920), .b(n784), .O(n940));
  inv1   g0639(.a(n920), .O(n941));
  nor2   g0640(.a(n941), .b(n783), .O(n942));
  nor2   g0641(.a(n942), .b(n926), .O(n943));
  inv1   g0642(.a(n943), .O(n944));
  nor2   g0643(.a(n944), .b(n940), .O(n945));
  inv1   g0644(.a(n410), .O(n946));
  nor2   g0645(.a(n930), .b(n946), .O(n947));
  inv1   g0646(.a(G129), .O(n948));
  nor2   g0647(.a(n935), .b(n948), .O(n949));
  nor2   g0648(.a(n949), .b(n947), .O(n950));
  inv1   g0649(.a(n950), .O(n951));
  nor2   g0650(.a(n951), .b(n945), .O(G838));
  inv1   g0651(.a(G4), .O(n953));
  nor2   g0652(.a(n669), .b(n666), .O(n954));
  inv1   g0653(.a(n954), .O(n955));
  nor2   g0654(.a(n955), .b(n953), .O(n956));
  nor2   g0655(.a(n954), .b(G4), .O(n957));
  nor2   g0656(.a(n957), .b(n956), .O(n958));
  inv1   g0657(.a(n958), .O(n959));
  nor2   g0658(.a(n959), .b(n926), .O(n960));
  inv1   g0659(.a(n561), .O(n961));
  nor2   g0660(.a(n930), .b(n961), .O(n962));
  inv1   g0661(.a(G117), .O(n963));
  nor2   g0662(.a(n935), .b(n963), .O(n964));
  nor2   g0663(.a(n964), .b(n962), .O(n965));
  inv1   g0664(.a(n965), .O(n966));
  nor2   g0665(.a(n966), .b(n960), .O(G861));
  nor2   g0666(.a(n806), .b(n795), .O(n968));
  inv1   g0667(.a(n968), .O(n969));
  inv1   g0668(.a(n940), .O(n970));
  nor2   g0669(.a(n970), .b(n776), .O(n971));
  inv1   g0670(.a(n971), .O(n972));
  nor2   g0671(.a(n972), .b(n922), .O(n973));
  nor2   g0672(.a(n973), .b(n809), .O(n974));
  nor2   g0673(.a(n974), .b(n969), .O(n975));
  nor2   g0674(.a(n975), .b(n806), .O(n976));
  nor2   g0675(.a(n976), .b(n805), .O(n977));
  nor2   g0676(.a(n977), .b(n802), .O(n978));
  nor2   g0677(.a(n978), .b(n766), .O(n979));
  nor2   g0678(.a(n979), .b(n915), .O(n980));
  inv1   g0679(.a(n980), .O(n981));
  nor2   g0680(.a(n743), .b(n739), .O(n982));
  nor2   g0681(.a(n982), .b(n745), .O(n983));
  nor2   g0682(.a(n983), .b(n981), .O(n984));
  nor2   g0683(.a(n980), .b(n743), .O(n985));
  nor2   g0684(.a(n985), .b(n984), .O(G623));
  inv1   g0685(.a(G4088), .O(n987));
  nor2   g0686(.a(n987), .b(G4087), .O(n988));
  inv1   g0687(.a(n988), .O(n989));
  nor2   g0688(.a(n989), .b(G861), .O(n990));
  nor2   g0689(.a(G4088), .b(G4087), .O(n991));
  inv1   g0690(.a(n991), .O(n992));
  nor2   g0691(.a(n992), .b(G822), .O(n993));
  nor2   g0692(.a(n987), .b(G61), .O(n994));
  inv1   g0693(.a(G4087), .O(n995));
  nor2   g0694(.a(G4088), .b(G11), .O(n996));
  nor2   g0695(.a(n996), .b(n995), .O(n997));
  inv1   g0696(.a(n997), .O(n998));
  nor2   g0697(.a(n998), .b(n994), .O(n999));
  nor2   g0698(.a(n999), .b(n993), .O(n1000));
  inv1   g0699(.a(n1000), .O(n1001));
  nor2   g0700(.a(n1001), .b(n990), .O(n1002));
  inv1   g0701(.a(n1002), .O(G722));
  inv1   g0702(.a(n976), .O(n1004));
  nor2   g0703(.a(n1004), .b(n804), .O(n1005));
  nor2   g0704(.a(n977), .b(n926), .O(n1006));
  inv1   g0705(.a(n1006), .O(n1007));
  nor2   g0706(.a(n1007), .b(n1005), .O(n1008));
  inv1   g0707(.a(n423), .O(n1009));
  nor2   g0708(.a(n930), .b(n1009), .O(n1010));
  inv1   g0709(.a(G52), .O(n1011));
  nor2   g0710(.a(n935), .b(n1011), .O(n1012));
  nor2   g0711(.a(n1012), .b(n1010), .O(n1013));
  inv1   g0712(.a(n1013), .O(n1014));
  nor2   g0713(.a(n1014), .b(n1008), .O(G832));
  inv1   g0714(.a(n974), .O(n1016));
  nor2   g0715(.a(n1016), .b(n968), .O(n1017));
  nor2   g0716(.a(n975), .b(n926), .O(n1018));
  inv1   g0717(.a(n1018), .O(n1019));
  nor2   g0718(.a(n1019), .b(n1017), .O(n1020));
  inv1   g0719(.a(n479), .O(n1021));
  nor2   g0720(.a(n930), .b(n1021), .O(n1022));
  inv1   g0721(.a(G130), .O(n1023));
  nor2   g0722(.a(n935), .b(n1023), .O(n1024));
  nor2   g0723(.a(n1024), .b(n1022), .O(n1025));
  inv1   g0724(.a(n1025), .O(n1026));
  nor2   g0725(.a(n1026), .b(n1020), .O(G834));
  nor2   g0726(.a(n782), .b(n776), .O(n1028));
  inv1   g0727(.a(n782), .O(n1029));
  nor2   g0728(.a(n1029), .b(n775), .O(n1030));
  nor2   g0729(.a(n1030), .b(n1028), .O(n1031));
  inv1   g0730(.a(n1031), .O(n1032));
  nor2   g0731(.a(n1032), .b(n940), .O(n1033));
  nor2   g0732(.a(n971), .b(n926), .O(n1034));
  inv1   g0733(.a(n1034), .O(n1035));
  nor2   g0734(.a(n1035), .b(n1033), .O(n1036));
  inv1   g0735(.a(n397), .O(n1037));
  nor2   g0736(.a(n930), .b(n1037), .O(n1038));
  inv1   g0737(.a(G119), .O(n1039));
  nor2   g0738(.a(n935), .b(n1039), .O(n1040));
  nor2   g0739(.a(n1040), .b(n1038), .O(n1041));
  inv1   g0740(.a(n1041), .O(n1042));
  nor2   g0741(.a(n1042), .b(n1036), .O(G836));
  inv1   g0742(.a(G4089), .O(n1044));
  nor2   g0743(.a(G4090), .b(n1044), .O(n1045));
  inv1   g0744(.a(n1045), .O(n1046));
  nor2   g0745(.a(n1046), .b(G861), .O(n1047));
  nor2   g0746(.a(G4090), .b(G4089), .O(n1048));
  inv1   g0747(.a(n1048), .O(n1049));
  nor2   g0748(.a(n1049), .b(G822), .O(n1050));
  nor2   g0749(.a(n1044), .b(G61), .O(n1051));
  inv1   g0750(.a(G4090), .O(n1052));
  nor2   g0751(.a(G4089), .b(G11), .O(n1053));
  nor2   g0752(.a(n1053), .b(n1052), .O(n1054));
  inv1   g0753(.a(n1054), .O(n1055));
  nor2   g0754(.a(n1055), .b(n1051), .O(n1056));
  nor2   g0755(.a(n1056), .b(n1050), .O(n1057));
  inv1   g0756(.a(n1057), .O(n1058));
  nor2   g0757(.a(n1058), .b(n1047), .O(n1059));
  inv1   g0758(.a(n1059), .O(G859));
  nor2   g0759(.a(n956), .b(n669), .O(n1061));
  nor2   g0760(.a(n1061), .b(n649), .O(n1062));
  nor2   g0761(.a(n1062), .b(n645), .O(n1063));
  nor2   g0762(.a(n1063), .b(n658), .O(n1064));
  nor2   g0763(.a(n1064), .b(n891), .O(n1065));
  nor2   g0764(.a(n1065), .b(n678), .O(n1066));
  nor2   g0765(.a(n1066), .b(n674), .O(n1067));
  nor2   g0766(.a(n1067), .b(n640), .O(n1068));
  inv1   g0767(.a(n1067), .O(n1069));
  nor2   g0768(.a(n1069), .b(n639), .O(n1070));
  nor2   g0769(.a(n1070), .b(n1068), .O(n1071));
  inv1   g0770(.a(n1071), .O(n1072));
  nor2   g0771(.a(n1072), .b(n926), .O(n1073));
  inv1   g0772(.a(n592), .O(n1074));
  nor2   g0773(.a(n930), .b(n1074), .O(n1075));
  inv1   g0774(.a(G122), .O(n1076));
  nor2   g0775(.a(n935), .b(n1076), .O(n1077));
  nor2   g0776(.a(n1077), .b(n1075), .O(n1078));
  inv1   g0777(.a(n1078), .O(n1079));
  nor2   g0778(.a(n1079), .b(n1073), .O(G871));
  inv1   g0779(.a(n1065), .O(n1081));
  nor2   g0780(.a(n1081), .b(n677), .O(n1082));
  nor2   g0781(.a(n1082), .b(n1066), .O(n1083));
  inv1   g0782(.a(n1083), .O(n1084));
  nor2   g0783(.a(n1084), .b(n926), .O(n1085));
  inv1   g0784(.a(n576), .O(n1086));
  nor2   g0785(.a(n930), .b(n1086), .O(n1087));
  inv1   g0786(.a(G128), .O(n1088));
  nor2   g0787(.a(n935), .b(n1088), .O(n1089));
  nor2   g0788(.a(n1089), .b(n1087), .O(n1090));
  inv1   g0789(.a(n1090), .O(n1091));
  nor2   g0790(.a(n1091), .b(n1085), .O(G873));
  inv1   g0791(.a(n1063), .O(n1093));
  nor2   g0792(.a(n1093), .b(n657), .O(n1094));
  nor2   g0793(.a(n1094), .b(n1064), .O(n1095));
  inv1   g0794(.a(n1095), .O(n1096));
  nor2   g0795(.a(n1096), .b(n926), .O(n1097));
  inv1   g0796(.a(n499), .O(n1098));
  nor2   g0797(.a(n930), .b(n1098), .O(n1099));
  inv1   g0798(.a(G127), .O(n1100));
  nor2   g0799(.a(n935), .b(n1100), .O(n1101));
  nor2   g0800(.a(n1101), .b(n1099), .O(n1102));
  inv1   g0801(.a(n1102), .O(n1103));
  nor2   g0802(.a(n1103), .b(n1097), .O(G875));
  inv1   g0803(.a(n1061), .O(n1105));
  nor2   g0804(.a(n1105), .b(n648), .O(n1106));
  nor2   g0805(.a(n1062), .b(n926), .O(n1107));
  inv1   g0806(.a(n1107), .O(n1108));
  nor2   g0807(.a(n1108), .b(n1106), .O(n1109));
  inv1   g0808(.a(n528), .O(n1110));
  nor2   g0809(.a(n930), .b(n1110), .O(n1111));
  inv1   g0810(.a(G126), .O(n1112));
  nor2   g0811(.a(n935), .b(n1112), .O(n1113));
  nor2   g0812(.a(n1113), .b(n1111), .O(n1114));
  inv1   g0813(.a(n1114), .O(n1115));
  nor2   g0814(.a(n1115), .b(n1109), .O(G877));
  inv1   g0815(.a(n983), .O(n1117));
  nor2   g0816(.a(n1117), .b(n759), .O(n1118));
  nor2   g0817(.a(n983), .b(n761), .O(n1119));
  nor2   g0818(.a(n1119), .b(n1118), .O(n1120));
  inv1   g0819(.a(n1120), .O(n1121));
  nor2   g0820(.a(n801), .b(n793), .O(n1122));
  nor2   g0821(.a(n794), .b(G331), .O(n1123));
  nor2   g0822(.a(n1123), .b(n1122), .O(n1124));
  nor2   g0823(.a(n1124), .b(n1121), .O(n1125));
  inv1   g0824(.a(n1124), .O(n1126));
  nor2   g0825(.a(n1126), .b(n1120), .O(n1127));
  nor2   g0826(.a(n1127), .b(n1125), .O(n1128));
  inv1   g0827(.a(n1128), .O(n1129));
  nor2   g0828(.a(G372), .b(n737), .O(n1130));
  nor2   g0829(.a(G369), .b(G332), .O(n1131));
  nor2   g0830(.a(n1131), .b(n1130), .O(n1132));
  nor2   g0831(.a(n1132), .b(n773), .O(n1133));
  inv1   g0832(.a(n1132), .O(n1134));
  nor2   g0833(.a(n1134), .b(n771), .O(n1135));
  nor2   g0834(.a(n1135), .b(n1133), .O(n1136));
  inv1   g0835(.a(n1136), .O(n1137));
  nor2   g0836(.a(n779), .b(n750), .O(n1138));
  nor2   g0837(.a(n780), .b(n752), .O(n1139));
  nor2   g0838(.a(n1139), .b(n1138), .O(n1140));
  nor2   g0839(.a(n1140), .b(n788), .O(n1141));
  inv1   g0840(.a(n1140), .O(n1142));
  nor2   g0841(.a(n1142), .b(n787), .O(n1143));
  nor2   g0842(.a(n1143), .b(n1141), .O(n1144));
  nor2   g0843(.a(n1144), .b(n1137), .O(n1145));
  inv1   g0844(.a(n1144), .O(n1146));
  nor2   g0845(.a(n1146), .b(n1136), .O(n1147));
  nor2   g0846(.a(n1147), .b(n1145), .O(n1148));
  inv1   g0847(.a(n1148), .O(n1149));
  nor2   g0848(.a(n1149), .b(n1129), .O(n1150));
  nor2   g0849(.a(n1148), .b(n1128), .O(n1151));
  nor2   g0850(.a(n1151), .b(n1150), .O(G998));
  nor2   g0851(.a(n664), .b(n653), .O(n1153));
  nor2   g0852(.a(n665), .b(n655), .O(n1154));
  nor2   g0853(.a(n1154), .b(n1153), .O(n1155));
  nor2   g0854(.a(n1155), .b(n637), .O(n1156));
  inv1   g0855(.a(n1155), .O(n1157));
  nor2   g0856(.a(n1157), .b(n635), .O(n1158));
  nor2   g0857(.a(n1158), .b(n1156), .O(n1159));
  inv1   g0858(.a(n1159), .O(n1160));
  nor2   g0859(.a(n697), .b(n688), .O(n1161));
  nor2   g0860(.a(n698), .b(n690), .O(n1162));
  nor2   g0861(.a(n1162), .b(n1161), .O(n1163));
  nor2   g0862(.a(n1163), .b(n705), .O(n1164));
  inv1   g0863(.a(n1163), .O(n1165));
  nor2   g0864(.a(n1165), .b(n703), .O(n1166));
  nor2   g0865(.a(n1166), .b(n1164), .O(n1167));
  inv1   g0866(.a(n1167), .O(n1168));
  nor2   g0867(.a(n673), .b(n644), .O(n1169));
  nor2   g0868(.a(n675), .b(n646), .O(n1170));
  nor2   g0869(.a(n1170), .b(n1169), .O(n1171));
  nor2   g0870(.a(n1171), .b(n720), .O(n1172));
  inv1   g0871(.a(n1171), .O(n1173));
  nor2   g0872(.a(n1173), .b(n718), .O(n1174));
  nor2   g0873(.a(n1174), .b(n1172), .O(n1175));
  inv1   g0874(.a(n1175), .O(n1176));
  nor2   g0875(.a(n1176), .b(n1168), .O(n1177));
  nor2   g0876(.a(n1175), .b(n1167), .O(n1178));
  nor2   g0877(.a(n1178), .b(n1177), .O(n1179));
  inv1   g0878(.a(n1179), .O(n1180));
  nor2   g0879(.a(n633), .b(G292), .O(n1181));
  nor2   g0880(.a(G335), .b(G289), .O(n1182));
  nor2   g0881(.a(n1182), .b(n1181), .O(n1183));
  nor2   g0882(.a(n1183), .b(n1180), .O(n1184));
  inv1   g0883(.a(n1183), .O(n1185));
  nor2   g0884(.a(n1185), .b(n1179), .O(n1186));
  nor2   g0885(.a(n1186), .b(n1184), .O(n1187));
  inv1   g0886(.a(n1187), .O(n1188));
  nor2   g0887(.a(n1188), .b(n1160), .O(n1189));
  nor2   g0888(.a(n1187), .b(n1159), .O(n1190));
  nor2   g0889(.a(n1190), .b(n1189), .O(n1191));
  inv1   g0890(.a(n1191), .O(G1000));
  inv1   g0891(.a(n898), .O(n1193));
  nor2   g0892(.a(n724), .b(n699), .O(n1194));
  inv1   g0893(.a(n1194), .O(n1195));
  nor2   g0894(.a(n1068), .b(n636), .O(n1196));
  nor2   g0895(.a(n1196), .b(n1195), .O(n1197));
  inv1   g0896(.a(n1197), .O(n1198));
  nor2   g0897(.a(n1198), .b(n708), .O(n1199));
  nor2   g0898(.a(n1199), .b(n1193), .O(n1200));
  inv1   g0899(.a(n1200), .O(n1201));
  nor2   g0900(.a(n1201), .b(n693), .O(n1202));
  nor2   g0901(.a(n1202), .b(n691), .O(n1203));
  inv1   g0902(.a(n1203), .O(n1204));
  nor2   g0903(.a(n1204), .b(n723), .O(n1205));
  nor2   g0904(.a(n1203), .b(n722), .O(n1206));
  nor2   g0905(.a(n1206), .b(n1205), .O(n1207));
  nor2   g0906(.a(n1200), .b(n692), .O(n1208));
  nor2   g0907(.a(n1208), .b(n1202), .O(n1209));
  inv1   g0908(.a(n1209), .O(n1210));
  nor2   g0909(.a(n1197), .b(n728), .O(n1211));
  nor2   g0910(.a(n1211), .b(n1199), .O(n1212));
  inv1   g0911(.a(n1196), .O(n1213));
  nor2   g0912(.a(n1213), .b(n1194), .O(n1214));
  nor2   g0913(.a(n1214), .b(n1197), .O(n1215));
  nor2   g0914(.a(n666), .b(n648), .O(n1216));
  inv1   g0915(.a(n666), .O(n1217));
  nor2   g0916(.a(n1217), .b(n649), .O(n1218));
  nor2   g0917(.a(n1218), .b(n1216), .O(n1219));
  inv1   g0918(.a(n1219), .O(n1220));
  nor2   g0919(.a(n1220), .b(n958), .O(n1221));
  inv1   g0920(.a(n1221), .O(n1222));
  nor2   g0921(.a(n1222), .b(n1095), .O(n1223));
  inv1   g0922(.a(n1223), .O(n1224));
  nor2   g0923(.a(n1224), .b(n1083), .O(n1225));
  inv1   g0924(.a(n1225), .O(n1226));
  nor2   g0925(.a(n1226), .b(n1071), .O(n1227));
  inv1   g0926(.a(n1227), .O(n1228));
  nor2   g0927(.a(n1228), .b(n1215), .O(n1229));
  inv1   g0928(.a(n1229), .O(n1230));
  nor2   g0929(.a(n1230), .b(n1212), .O(n1231));
  inv1   g0930(.a(n1231), .O(n1232));
  nor2   g0931(.a(n1232), .b(n1210), .O(n1233));
  inv1   g0932(.a(n1233), .O(n1234));
  nor2   g0933(.a(n1234), .b(n1207), .O(G575));
  nor2   g0934(.a(n981), .b(n740), .O(n1236));
  nor2   g0935(.a(n980), .b(n739), .O(n1237));
  nor2   g0936(.a(n1237), .b(n1236), .O(n1238));
  inv1   g0937(.a(n1238), .O(n1239));
  inv1   g0938(.a(G623), .O(n1240));
  inv1   g0939(.a(n973), .O(n1241));
  nor2   g0940(.a(n969), .b(n805), .O(n1242));
  inv1   g0941(.a(n1242), .O(n1243));
  nor2   g0942(.a(n1243), .b(n766), .O(n1244));
  inv1   g0943(.a(n1244), .O(n1245));
  nor2   g0944(.a(n1245), .b(n1241), .O(n1246));
  inv1   g0945(.a(n1246), .O(n1247));
  nor2   g0946(.a(n1247), .b(n1240), .O(n1248));
  inv1   g0947(.a(n1248), .O(n1249));
  nor2   g0948(.a(n1249), .b(n1239), .O(G585));
  inv1   g0949(.a(G137), .O(n1251));
  inv1   g0950(.a(G1689), .O(n1252));
  nor2   g0951(.a(G1690), .b(n1252), .O(n1253));
  inv1   g0952(.a(n1253), .O(n1254));
  nor2   g0953(.a(n1254), .b(G861), .O(n1255));
  nor2   g0954(.a(G1690), .b(G1689), .O(n1256));
  inv1   g0955(.a(n1256), .O(n1257));
  nor2   g0956(.a(n1257), .b(G822), .O(n1258));
  nor2   g0957(.a(n1252), .b(G185), .O(n1259));
  inv1   g0958(.a(G1690), .O(n1260));
  nor2   g0959(.a(G1689), .b(G182), .O(n1261));
  nor2   g0960(.a(n1261), .b(n1260), .O(n1262));
  inv1   g0961(.a(n1262), .O(n1263));
  nor2   g0962(.a(n1263), .b(n1259), .O(n1264));
  nor2   g0963(.a(n1264), .b(n1258), .O(n1265));
  inv1   g0964(.a(n1265), .O(n1266));
  nor2   g0965(.a(n1266), .b(n1255), .O(n1267));
  nor2   g0966(.a(n1267), .b(n1251), .O(G661));
  inv1   g0967(.a(G1691), .O(n1269));
  nor2   g0968(.a(G1694), .b(n1269), .O(n1270));
  inv1   g0969(.a(n1270), .O(n1271));
  nor2   g0970(.a(n1271), .b(G861), .O(n1272));
  nor2   g0971(.a(G1694), .b(G1691), .O(n1273));
  inv1   g0972(.a(n1273), .O(n1274));
  nor2   g0973(.a(n1274), .b(G822), .O(n1275));
  nor2   g0974(.a(n1269), .b(G185), .O(n1276));
  inv1   g0975(.a(G1694), .O(n1277));
  nor2   g0976(.a(G1691), .b(G182), .O(n1278));
  nor2   g0977(.a(n1278), .b(n1277), .O(n1279));
  inv1   g0978(.a(n1279), .O(n1280));
  nor2   g0979(.a(n1280), .b(n1276), .O(n1281));
  nor2   g0980(.a(n1281), .b(n1275), .O(n1282));
  inv1   g0981(.a(n1282), .O(n1283));
  nor2   g0982(.a(n1283), .b(n1272), .O(n1284));
  nor2   g0983(.a(n1284), .b(n1251), .O(G693));
  nor2   g0984(.a(G871), .b(n989), .O(n1286));
  nor2   g0985(.a(G832), .b(n992), .O(n1287));
  nor2   g0986(.a(n987), .b(G37), .O(n1288));
  nor2   g0987(.a(G4088), .b(G43), .O(n1289));
  nor2   g0988(.a(n1289), .b(n995), .O(n1290));
  inv1   g0989(.a(n1290), .O(n1291));
  nor2   g0990(.a(n1291), .b(n1288), .O(n1292));
  nor2   g0991(.a(n1292), .b(n1287), .O(n1293));
  inv1   g0992(.a(n1293), .O(n1294));
  nor2   g0993(.a(n1294), .b(n1286), .O(n1295));
  inv1   g0994(.a(n1295), .O(G747));
  nor2   g0995(.a(G873), .b(n989), .O(n1297));
  nor2   g0996(.a(G834), .b(n992), .O(n1298));
  nor2   g0997(.a(n987), .b(G20), .O(n1299));
  nor2   g0998(.a(G4088), .b(G76), .O(n1300));
  nor2   g0999(.a(n1300), .b(n995), .O(n1301));
  inv1   g1000(.a(n1301), .O(n1302));
  nor2   g1001(.a(n1302), .b(n1299), .O(n1303));
  nor2   g1002(.a(n1303), .b(n1298), .O(n1304));
  inv1   g1003(.a(n1304), .O(n1305));
  nor2   g1004(.a(n1305), .b(n1297), .O(n1306));
  inv1   g1005(.a(n1306), .O(G752));
  nor2   g1006(.a(G875), .b(n989), .O(n1308));
  nor2   g1007(.a(G836), .b(n992), .O(n1309));
  nor2   g1008(.a(n987), .b(G17), .O(n1310));
  nor2   g1009(.a(G4088), .b(G73), .O(n1311));
  nor2   g1010(.a(n1311), .b(n995), .O(n1312));
  inv1   g1011(.a(n1312), .O(n1313));
  nor2   g1012(.a(n1313), .b(n1310), .O(n1314));
  nor2   g1013(.a(n1314), .b(n1309), .O(n1315));
  inv1   g1014(.a(n1315), .O(n1316));
  nor2   g1015(.a(n1316), .b(n1308), .O(n1317));
  inv1   g1016(.a(n1317), .O(G757));
  nor2   g1017(.a(G877), .b(n989), .O(n1319));
  nor2   g1018(.a(n992), .b(G838), .O(n1320));
  nor2   g1019(.a(n987), .b(G70), .O(n1321));
  nor2   g1020(.a(G4088), .b(G67), .O(n1322));
  nor2   g1021(.a(n1322), .b(n995), .O(n1323));
  inv1   g1022(.a(n1323), .O(n1324));
  nor2   g1023(.a(n1324), .b(n1321), .O(n1325));
  nor2   g1024(.a(n1325), .b(n1320), .O(n1326));
  inv1   g1025(.a(n1326), .O(n1327));
  nor2   g1026(.a(n1327), .b(n1319), .O(n1328));
  inv1   g1027(.a(n1328), .O(G762));
  nor2   g1028(.a(G871), .b(n1046), .O(n1330));
  nor2   g1029(.a(n1049), .b(G832), .O(n1331));
  nor2   g1030(.a(n1044), .b(G37), .O(n1332));
  nor2   g1031(.a(G4089), .b(G43), .O(n1333));
  nor2   g1032(.a(n1333), .b(n1052), .O(n1334));
  inv1   g1033(.a(n1334), .O(n1335));
  nor2   g1034(.a(n1335), .b(n1332), .O(n1336));
  nor2   g1035(.a(n1336), .b(n1331), .O(n1337));
  inv1   g1036(.a(n1337), .O(n1338));
  nor2   g1037(.a(n1338), .b(n1330), .O(n1339));
  inv1   g1038(.a(n1339), .O(G787));
  nor2   g1039(.a(G873), .b(n1046), .O(n1341));
  nor2   g1040(.a(n1049), .b(G834), .O(n1342));
  nor2   g1041(.a(n1044), .b(G20), .O(n1343));
  nor2   g1042(.a(G4089), .b(G76), .O(n1344));
  nor2   g1043(.a(n1344), .b(n1052), .O(n1345));
  inv1   g1044(.a(n1345), .O(n1346));
  nor2   g1045(.a(n1346), .b(n1343), .O(n1347));
  nor2   g1046(.a(n1347), .b(n1342), .O(n1348));
  inv1   g1047(.a(n1348), .O(n1349));
  nor2   g1048(.a(n1349), .b(n1341), .O(n1350));
  inv1   g1049(.a(n1350), .O(G792));
  nor2   g1050(.a(G875), .b(n1046), .O(n1352));
  nor2   g1051(.a(n1049), .b(G836), .O(n1353));
  nor2   g1052(.a(n1044), .b(G17), .O(n1354));
  nor2   g1053(.a(G4089), .b(G73), .O(n1355));
  nor2   g1054(.a(n1355), .b(n1052), .O(n1356));
  inv1   g1055(.a(n1356), .O(n1357));
  nor2   g1056(.a(n1357), .b(n1354), .O(n1358));
  nor2   g1057(.a(n1358), .b(n1353), .O(n1359));
  inv1   g1058(.a(n1359), .O(n1360));
  nor2   g1059(.a(n1360), .b(n1352), .O(n1361));
  inv1   g1060(.a(n1361), .O(G797));
  nor2   g1061(.a(G877), .b(n1046), .O(n1363));
  nor2   g1062(.a(n1049), .b(G838), .O(n1364));
  nor2   g1063(.a(n1044), .b(G70), .O(n1365));
  nor2   g1064(.a(G4089), .b(G67), .O(n1366));
  nor2   g1065(.a(n1366), .b(n1052), .O(n1367));
  inv1   g1066(.a(n1367), .O(n1368));
  nor2   g1067(.a(n1368), .b(n1365), .O(n1369));
  nor2   g1068(.a(n1369), .b(n1364), .O(n1370));
  inv1   g1069(.a(n1370), .O(n1371));
  nor2   g1070(.a(n1371), .b(n1363), .O(n1372));
  inv1   g1071(.a(n1372), .O(G802));
  nor2   g1072(.a(n1254), .b(G871), .O(n1374));
  nor2   g1073(.a(n1257), .b(G832), .O(n1375));
  nor2   g1074(.a(n1252), .b(G170), .O(n1376));
  nor2   g1075(.a(G1689), .b(G200), .O(n1377));
  nor2   g1076(.a(n1377), .b(n1260), .O(n1378));
  inv1   g1077(.a(n1378), .O(n1379));
  nor2   g1078(.a(n1379), .b(n1376), .O(n1380));
  nor2   g1079(.a(n1380), .b(n1375), .O(n1381));
  inv1   g1080(.a(n1381), .O(n1382));
  nor2   g1081(.a(n1382), .b(n1374), .O(n1383));
  nor2   g1082(.a(n1383), .b(n1251), .O(G642));
  nor2   g1083(.a(n1254), .b(G877), .O(n1385));
  nor2   g1084(.a(n1257), .b(G838), .O(n1386));
  nor2   g1085(.a(n1252), .b(G158), .O(n1387));
  nor2   g1086(.a(G1689), .b(G188), .O(n1388));
  nor2   g1087(.a(n1388), .b(n1260), .O(n1389));
  inv1   g1088(.a(n1389), .O(n1390));
  nor2   g1089(.a(n1390), .b(n1387), .O(n1391));
  nor2   g1090(.a(n1391), .b(n1386), .O(n1392));
  inv1   g1091(.a(n1392), .O(n1393));
  nor2   g1092(.a(n1393), .b(n1385), .O(n1394));
  nor2   g1093(.a(n1394), .b(n1251), .O(G664));
  nor2   g1094(.a(n1254), .b(G875), .O(n1396));
  nor2   g1095(.a(n1257), .b(G836), .O(n1397));
  nor2   g1096(.a(n1252), .b(G152), .O(n1398));
  nor2   g1097(.a(G1689), .b(G155), .O(n1399));
  nor2   g1098(.a(n1399), .b(n1260), .O(n1400));
  inv1   g1099(.a(n1400), .O(n1401));
  nor2   g1100(.a(n1401), .b(n1398), .O(n1402));
  nor2   g1101(.a(n1402), .b(n1397), .O(n1403));
  inv1   g1102(.a(n1403), .O(n1404));
  nor2   g1103(.a(n1404), .b(n1396), .O(n1405));
  nor2   g1104(.a(n1405), .b(n1251), .O(G667));
  nor2   g1105(.a(n1254), .b(G873), .O(n1407));
  nor2   g1106(.a(n1257), .b(G834), .O(n1408));
  nor2   g1107(.a(n1252), .b(G146), .O(n1409));
  nor2   g1108(.a(G1689), .b(G149), .O(n1410));
  nor2   g1109(.a(n1410), .b(n1260), .O(n1411));
  inv1   g1110(.a(n1411), .O(n1412));
  nor2   g1111(.a(n1412), .b(n1409), .O(n1413));
  nor2   g1112(.a(n1413), .b(n1408), .O(n1414));
  inv1   g1113(.a(n1414), .O(n1415));
  nor2   g1114(.a(n1415), .b(n1407), .O(n1416));
  nor2   g1115(.a(n1416), .b(n1251), .O(G670));
  nor2   g1116(.a(n1271), .b(G871), .O(n1418));
  nor2   g1117(.a(n1274), .b(G832), .O(n1419));
  nor2   g1118(.a(n1269), .b(G170), .O(n1420));
  nor2   g1119(.a(G1691), .b(G200), .O(n1421));
  nor2   g1120(.a(n1421), .b(n1277), .O(n1422));
  inv1   g1121(.a(n1422), .O(n1423));
  nor2   g1122(.a(n1423), .b(n1420), .O(n1424));
  nor2   g1123(.a(n1424), .b(n1419), .O(n1425));
  inv1   g1124(.a(n1425), .O(n1426));
  nor2   g1125(.a(n1426), .b(n1418), .O(n1427));
  nor2   g1126(.a(n1427), .b(n1251), .O(G676));
  nor2   g1127(.a(n1271), .b(G877), .O(n1429));
  nor2   g1128(.a(n1274), .b(G838), .O(n1430));
  nor2   g1129(.a(n1269), .b(G158), .O(n1431));
  nor2   g1130(.a(G1691), .b(G188), .O(n1432));
  nor2   g1131(.a(n1432), .b(n1277), .O(n1433));
  inv1   g1132(.a(n1433), .O(n1434));
  nor2   g1133(.a(n1434), .b(n1431), .O(n1435));
  nor2   g1134(.a(n1435), .b(n1430), .O(n1436));
  inv1   g1135(.a(n1436), .O(n1437));
  nor2   g1136(.a(n1437), .b(n1429), .O(n1438));
  nor2   g1137(.a(n1438), .b(n1251), .O(G696));
  nor2   g1138(.a(n1271), .b(G875), .O(n1440));
  nor2   g1139(.a(n1274), .b(G836), .O(n1441));
  nor2   g1140(.a(n1269), .b(G152), .O(n1442));
  nor2   g1141(.a(G1691), .b(G155), .O(n1443));
  nor2   g1142(.a(n1443), .b(n1277), .O(n1444));
  inv1   g1143(.a(n1444), .O(n1445));
  nor2   g1144(.a(n1445), .b(n1442), .O(n1446));
  nor2   g1145(.a(n1446), .b(n1441), .O(n1447));
  inv1   g1146(.a(n1447), .O(n1448));
  nor2   g1147(.a(n1448), .b(n1440), .O(n1449));
  nor2   g1148(.a(n1449), .b(n1251), .O(G699));
  nor2   g1149(.a(n1271), .b(G873), .O(n1451));
  nor2   g1150(.a(n1274), .b(G834), .O(n1452));
  nor2   g1151(.a(n1269), .b(G146), .O(n1453));
  nor2   g1152(.a(G1691), .b(G149), .O(n1454));
  nor2   g1153(.a(n1454), .b(n1277), .O(n1455));
  inv1   g1154(.a(n1455), .O(n1456));
  nor2   g1155(.a(n1456), .b(n1453), .O(n1457));
  nor2   g1156(.a(n1457), .b(n1452), .O(n1458));
  inv1   g1157(.a(n1458), .O(n1459));
  nor2   g1158(.a(n1459), .b(n1451), .O(n1460));
  nor2   g1159(.a(n1460), .b(n1251), .O(G702));
  inv1   g1160(.a(G3724), .O(n1462));
  nor2   g1161(.a(G623), .b(n1462), .O(n1463));
  inv1   g1162(.a(G3717), .O(n1464));
  inv1   g1163(.a(G123), .O(n1465));
  nor2   g1164(.a(G3724), .b(n1465), .O(n1466));
  nor2   g1165(.a(n1466), .b(n1464), .O(n1467));
  inv1   g1166(.a(n1467), .O(n1468));
  nor2   g1167(.a(n1468), .b(n1463), .O(n1469));
  inv1   g1168(.a(G135), .O(n1470));
  inv1   g1169(.a(G4115), .O(n1471));
  nor2   g1170(.a(n1471), .b(n1470), .O(n1472));
  inv1   g1171(.a(G132), .O(n1473));
  nor2   g1172(.a(n743), .b(n1473), .O(n1474));
  nor2   g1173(.a(n744), .b(G132), .O(n1475));
  nor2   g1174(.a(n1475), .b(n1474), .O(n1476));
  nor2   g1175(.a(n1476), .b(n1462), .O(n1477));
  nor2   g1176(.a(n471), .b(G3724), .O(n1478));
  nor2   g1177(.a(n1478), .b(G3717), .O(n1479));
  inv1   g1178(.a(n1479), .O(n1480));
  nor2   g1179(.a(n1480), .b(n1477), .O(n1481));
  nor2   g1180(.a(n1481), .b(n1472), .O(n1482));
  inv1   g1181(.a(n1482), .O(n1483));
  nor2   g1182(.a(n1483), .b(n1469), .O(G818));
  nor2   g1183(.a(n1236), .b(n1473), .O(n1485));
  inv1   g1184(.a(n1236), .O(n1486));
  nor2   g1185(.a(n1486), .b(G132), .O(n1487));
  nor2   g1186(.a(n1487), .b(n1485), .O(G813));
  nor2   g1187(.a(G623), .b(n926), .O(n1489));
  nor2   g1188(.a(n930), .b(n471), .O(n1490));
  nor2   g1189(.a(n935), .b(n1465), .O(n1491));
  nor2   g1190(.a(n1491), .b(n1490), .O(n1492));
  inv1   g1191(.a(n1492), .O(n1493));
  nor2   g1192(.a(n1493), .b(n1489), .O(G824));
  nor2   g1193(.a(n1238), .b(n926), .O(n1495));
  inv1   g1194(.a(n433), .O(n1496));
  nor2   g1195(.a(n930), .b(n1496), .O(n1497));
  inv1   g1196(.a(G121), .O(n1498));
  nor2   g1197(.a(n935), .b(n1498), .O(n1499));
  nor2   g1198(.a(n1499), .b(n1497), .O(n1500));
  inv1   g1199(.a(n1500), .O(n1501));
  nor2   g1200(.a(n1501), .b(n1495), .O(G826));
  inv1   g1201(.a(n978), .O(n1503));
  nor2   g1202(.a(n1503), .b(n755), .O(n1504));
  inv1   g1203(.a(n753), .O(n1505));
  nor2   g1204(.a(n764), .b(n1505), .O(n1506));
  nor2   g1205(.a(n763), .b(n753), .O(n1507));
  nor2   g1206(.a(n1507), .b(n1506), .O(n1508));
  inv1   g1207(.a(n1508), .O(n1509));
  nor2   g1208(.a(n1509), .b(n1504), .O(n1510));
  inv1   g1209(.a(n1504), .O(n1511));
  nor2   g1210(.a(n1511), .b(n763), .O(n1512));
  nor2   g1211(.a(n1512), .b(n926), .O(n1513));
  inv1   g1212(.a(n1513), .O(n1514));
  nor2   g1213(.a(n1514), .b(n1510), .O(n1515));
  inv1   g1214(.a(n448), .O(n1516));
  nor2   g1215(.a(n930), .b(n1516), .O(n1517));
  inv1   g1216(.a(G116), .O(n1518));
  nor2   g1217(.a(n935), .b(n1518), .O(n1519));
  nor2   g1218(.a(n1519), .b(n1517), .O(n1520));
  inv1   g1219(.a(n1520), .O(n1521));
  nor2   g1220(.a(n1521), .b(n1515), .O(G828));
  nor2   g1221(.a(n978), .b(n754), .O(n1523));
  nor2   g1222(.a(n1523), .b(n1504), .O(n1524));
  nor2   g1223(.a(n1524), .b(n926), .O(n1525));
  inv1   g1224(.a(n463), .O(n1526));
  nor2   g1225(.a(n930), .b(n1526), .O(n1527));
  inv1   g1226(.a(G112), .O(n1528));
  nor2   g1227(.a(n935), .b(n1528), .O(n1529));
  nor2   g1228(.a(n1529), .b(n1527), .O(n1530));
  inv1   g1229(.a(n1530), .O(n1531));
  nor2   g1230(.a(n1531), .b(n1525), .O(G830));
  inv1   g1231(.a(G601), .O(n1533));
  nor2   g1232(.a(G851), .b(G848), .O(n1534));
  inv1   g1233(.a(n1534), .O(n1535));
  nor2   g1234(.a(n1535), .b(n1533), .O(n1536));
  inv1   g1235(.a(n1536), .O(n1537));
  nor2   g1236(.a(n1537), .b(G847), .O(n1538));
  inv1   g1237(.a(n1538), .O(n1539));
  nor2   g1238(.a(n1539), .b(G1002), .O(n1540));
  inv1   g1239(.a(n1540), .O(n1541));
  nor2   g1240(.a(n1541), .b(G1004), .O(n1542));
  inv1   g1241(.a(n1542), .O(n1543));
  nor2   g1242(.a(n1543), .b(G998), .O(n1544));
  inv1   g1243(.a(n1544), .O(n1545));
  nor2   g1244(.a(n1545), .b(G1000), .O(G854));
  inv1   g1245(.a(n1207), .O(n1547));
  nor2   g1246(.a(n1547), .b(n926), .O(n1548));
  inv1   g1247(.a(n607), .O(n1549));
  nor2   g1248(.a(n930), .b(n1549), .O(n1550));
  inv1   g1249(.a(G115), .O(n1551));
  nor2   g1250(.a(n935), .b(n1551), .O(n1552));
  nor2   g1251(.a(n1552), .b(n1550), .O(n1553));
  inv1   g1252(.a(n1553), .O(n1554));
  nor2   g1253(.a(n1554), .b(n1548), .O(G863));
  nor2   g1254(.a(n1209), .b(n926), .O(n1556));
  inv1   g1255(.a(n515), .O(n1557));
  nor2   g1256(.a(n930), .b(n1557), .O(n1558));
  inv1   g1257(.a(G114), .O(n1559));
  nor2   g1258(.a(n935), .b(n1559), .O(n1560));
  nor2   g1259(.a(n1560), .b(n1558), .O(n1561));
  inv1   g1260(.a(n1561), .O(n1562));
  nor2   g1261(.a(n1562), .b(n1556), .O(G865));
  inv1   g1262(.a(n1212), .O(n1564));
  nor2   g1263(.a(n1564), .b(n926), .O(n1565));
  inv1   g1264(.a(n623), .O(n1566));
  nor2   g1265(.a(n930), .b(n1566), .O(n1567));
  inv1   g1266(.a(G53), .O(n1568));
  nor2   g1267(.a(n935), .b(n1568), .O(n1569));
  nor2   g1268(.a(n1569), .b(n1567), .O(n1570));
  inv1   g1269(.a(n1570), .O(n1571));
  nor2   g1270(.a(n1571), .b(n1565), .O(G867));
  inv1   g1271(.a(n1215), .O(n1573));
  nor2   g1272(.a(n1573), .b(n926), .O(n1574));
  inv1   g1273(.a(n548), .O(n1575));
  nor2   g1274(.a(n930), .b(n1575), .O(n1576));
  inv1   g1275(.a(G113), .O(n1577));
  nor2   g1276(.a(n935), .b(n1577), .O(n1578));
  nor2   g1277(.a(n1578), .b(n1576), .O(n1579));
  inv1   g1278(.a(n1579), .O(n1580));
  nor2   g1279(.a(n1580), .b(n1574), .O(G869));
  nor2   g1280(.a(G863), .b(n1046), .O(n1582));
  nor2   g1281(.a(G824), .b(n1049), .O(n1583));
  nor2   g1282(.a(n1044), .b(G106), .O(n1584));
  nor2   g1283(.a(G4089), .b(G109), .O(n1585));
  nor2   g1284(.a(n1585), .b(n1052), .O(n1586));
  inv1   g1285(.a(n1586), .O(n1587));
  nor2   g1286(.a(n1587), .b(n1584), .O(n1588));
  nor2   g1287(.a(n1588), .b(n1583), .O(n1589));
  inv1   g1288(.a(n1589), .O(n1590));
  nor2   g1289(.a(n1590), .b(n1582), .O(n1591));
  inv1   g1290(.a(n1591), .O(G712));
  nor2   g1291(.a(G863), .b(n989), .O(n1593));
  nor2   g1292(.a(G824), .b(n992), .O(n1594));
  nor2   g1293(.a(n987), .b(G106), .O(n1595));
  nor2   g1294(.a(G4088), .b(G109), .O(n1596));
  nor2   g1295(.a(n1596), .b(n995), .O(n1597));
  inv1   g1296(.a(n1597), .O(n1598));
  nor2   g1297(.a(n1598), .b(n1595), .O(n1599));
  nor2   g1298(.a(n1599), .b(n1594), .O(n1600));
  inv1   g1299(.a(n1600), .O(n1601));
  nor2   g1300(.a(n1601), .b(n1593), .O(n1602));
  inv1   g1301(.a(n1602), .O(G727));
  nor2   g1302(.a(G865), .b(n989), .O(n1604));
  nor2   g1303(.a(G826), .b(n992), .O(n1605));
  nor2   g1304(.a(n987), .b(G49), .O(n1606));
  nor2   g1305(.a(G4088), .b(G46), .O(n1607));
  nor2   g1306(.a(n1607), .b(n995), .O(n1608));
  inv1   g1307(.a(n1608), .O(n1609));
  nor2   g1308(.a(n1609), .b(n1606), .O(n1610));
  nor2   g1309(.a(n1610), .b(n1605), .O(n1611));
  inv1   g1310(.a(n1611), .O(n1612));
  nor2   g1311(.a(n1612), .b(n1604), .O(n1613));
  inv1   g1312(.a(n1613), .O(G732));
  nor2   g1313(.a(G867), .b(n989), .O(n1615));
  nor2   g1314(.a(G828), .b(n992), .O(n1616));
  nor2   g1315(.a(n987), .b(G103), .O(n1617));
  nor2   g1316(.a(G4088), .b(G100), .O(n1618));
  nor2   g1317(.a(n1618), .b(n995), .O(n1619));
  inv1   g1318(.a(n1619), .O(n1620));
  nor2   g1319(.a(n1620), .b(n1617), .O(n1621));
  nor2   g1320(.a(n1621), .b(n1616), .O(n1622));
  inv1   g1321(.a(n1622), .O(n1623));
  nor2   g1322(.a(n1623), .b(n1615), .O(n1624));
  inv1   g1323(.a(n1624), .O(G737));
  nor2   g1324(.a(G869), .b(n989), .O(n1626));
  nor2   g1325(.a(G830), .b(n992), .O(n1627));
  nor2   g1326(.a(n987), .b(G40), .O(n1628));
  nor2   g1327(.a(G4088), .b(G91), .O(n1629));
  nor2   g1328(.a(n1629), .b(n995), .O(n1630));
  inv1   g1329(.a(n1630), .O(n1631));
  nor2   g1330(.a(n1631), .b(n1628), .O(n1632));
  nor2   g1331(.a(n1632), .b(n1627), .O(n1633));
  inv1   g1332(.a(n1633), .O(n1634));
  nor2   g1333(.a(n1634), .b(n1626), .O(n1635));
  inv1   g1334(.a(n1635), .O(G742));
  nor2   g1335(.a(G865), .b(n1046), .O(n1637));
  nor2   g1336(.a(G826), .b(n1049), .O(n1638));
  nor2   g1337(.a(n1044), .b(G49), .O(n1639));
  nor2   g1338(.a(G4089), .b(G46), .O(n1640));
  nor2   g1339(.a(n1640), .b(n1052), .O(n1641));
  inv1   g1340(.a(n1641), .O(n1642));
  nor2   g1341(.a(n1642), .b(n1639), .O(n1643));
  nor2   g1342(.a(n1643), .b(n1638), .O(n1644));
  inv1   g1343(.a(n1644), .O(n1645));
  nor2   g1344(.a(n1645), .b(n1637), .O(n1646));
  inv1   g1345(.a(n1646), .O(G772));
  nor2   g1346(.a(G867), .b(n1046), .O(n1648));
  nor2   g1347(.a(G828), .b(n1049), .O(n1649));
  nor2   g1348(.a(n1044), .b(G103), .O(n1650));
  nor2   g1349(.a(G4089), .b(G100), .O(n1651));
  nor2   g1350(.a(n1651), .b(n1052), .O(n1652));
  inv1   g1351(.a(n1652), .O(n1653));
  nor2   g1352(.a(n1653), .b(n1650), .O(n1654));
  nor2   g1353(.a(n1654), .b(n1649), .O(n1655));
  inv1   g1354(.a(n1655), .O(n1656));
  nor2   g1355(.a(n1656), .b(n1648), .O(n1657));
  inv1   g1356(.a(n1657), .O(G777));
  nor2   g1357(.a(G869), .b(n1046), .O(n1659));
  nor2   g1358(.a(G830), .b(n1049), .O(n1660));
  nor2   g1359(.a(n1044), .b(G40), .O(n1661));
  nor2   g1360(.a(G4089), .b(G91), .O(n1662));
  nor2   g1361(.a(n1662), .b(n1052), .O(n1663));
  inv1   g1362(.a(n1663), .O(n1664));
  nor2   g1363(.a(n1664), .b(n1661), .O(n1665));
  nor2   g1364(.a(n1665), .b(n1660), .O(n1666));
  inv1   g1365(.a(n1666), .O(n1667));
  nor2   g1366(.a(n1667), .b(n1659), .O(n1668));
  inv1   g1367(.a(n1668), .O(G782));
  nor2   g1368(.a(G869), .b(n1254), .O(n1670));
  nor2   g1369(.a(G830), .b(n1257), .O(n1671));
  nor2   g1370(.a(n1252), .b(G173), .O(n1672));
  nor2   g1371(.a(G1689), .b(G203), .O(n1673));
  nor2   g1372(.a(n1673), .b(n1260), .O(n1674));
  inv1   g1373(.a(n1674), .O(n1675));
  nor2   g1374(.a(n1675), .b(n1672), .O(n1676));
  nor2   g1375(.a(n1676), .b(n1671), .O(n1677));
  inv1   g1376(.a(n1677), .O(n1678));
  nor2   g1377(.a(n1678), .b(n1670), .O(n1679));
  nor2   g1378(.a(n1679), .b(n1251), .O(G645));
  nor2   g1379(.a(G867), .b(n1254), .O(n1681));
  nor2   g1380(.a(G828), .b(n1257), .O(n1682));
  nor2   g1381(.a(n1252), .b(G167), .O(n1683));
  nor2   g1382(.a(G1689), .b(G197), .O(n1684));
  nor2   g1383(.a(n1684), .b(n1260), .O(n1685));
  inv1   g1384(.a(n1685), .O(n1686));
  nor2   g1385(.a(n1686), .b(n1683), .O(n1687));
  nor2   g1386(.a(n1687), .b(n1682), .O(n1688));
  inv1   g1387(.a(n1688), .O(n1689));
  nor2   g1388(.a(n1689), .b(n1681), .O(n1690));
  nor2   g1389(.a(n1690), .b(n1251), .O(G648));
  nor2   g1390(.a(G865), .b(n1254), .O(n1692));
  nor2   g1391(.a(G826), .b(n1257), .O(n1693));
  nor2   g1392(.a(n1252), .b(G164), .O(n1694));
  nor2   g1393(.a(G1689), .b(G194), .O(n1695));
  nor2   g1394(.a(n1695), .b(n1260), .O(n1696));
  inv1   g1395(.a(n1696), .O(n1697));
  nor2   g1396(.a(n1697), .b(n1694), .O(n1698));
  nor2   g1397(.a(n1698), .b(n1693), .O(n1699));
  inv1   g1398(.a(n1699), .O(n1700));
  nor2   g1399(.a(n1700), .b(n1692), .O(n1701));
  nor2   g1400(.a(n1701), .b(n1251), .O(G651));
  nor2   g1401(.a(G863), .b(n1254), .O(n1703));
  nor2   g1402(.a(G824), .b(n1257), .O(n1704));
  nor2   g1403(.a(n1252), .b(G161), .O(n1705));
  nor2   g1404(.a(G1689), .b(G191), .O(n1706));
  nor2   g1405(.a(n1706), .b(n1260), .O(n1707));
  inv1   g1406(.a(n1707), .O(n1708));
  nor2   g1407(.a(n1708), .b(n1705), .O(n1709));
  nor2   g1408(.a(n1709), .b(n1704), .O(n1710));
  inv1   g1409(.a(n1710), .O(n1711));
  nor2   g1410(.a(n1711), .b(n1703), .O(n1712));
  nor2   g1411(.a(n1712), .b(n1251), .O(G654));
  nor2   g1412(.a(G869), .b(n1271), .O(n1714));
  nor2   g1413(.a(G830), .b(n1274), .O(n1715));
  nor2   g1414(.a(n1269), .b(G173), .O(n1716));
  nor2   g1415(.a(G1691), .b(G203), .O(n1717));
  nor2   g1416(.a(n1717), .b(n1277), .O(n1718));
  inv1   g1417(.a(n1718), .O(n1719));
  nor2   g1418(.a(n1719), .b(n1716), .O(n1720));
  nor2   g1419(.a(n1720), .b(n1715), .O(n1721));
  inv1   g1420(.a(n1721), .O(n1722));
  nor2   g1421(.a(n1722), .b(n1714), .O(n1723));
  nor2   g1422(.a(n1723), .b(n1251), .O(G679));
  nor2   g1423(.a(G867), .b(n1271), .O(n1725));
  nor2   g1424(.a(G828), .b(n1274), .O(n1726));
  nor2   g1425(.a(n1269), .b(G167), .O(n1727));
  nor2   g1426(.a(G1691), .b(G197), .O(n1728));
  nor2   g1427(.a(n1728), .b(n1277), .O(n1729));
  inv1   g1428(.a(n1729), .O(n1730));
  nor2   g1429(.a(n1730), .b(n1727), .O(n1731));
  nor2   g1430(.a(n1731), .b(n1726), .O(n1732));
  inv1   g1431(.a(n1732), .O(n1733));
  nor2   g1432(.a(n1733), .b(n1725), .O(n1734));
  nor2   g1433(.a(n1734), .b(n1251), .O(G682));
  nor2   g1434(.a(G865), .b(n1271), .O(n1736));
  nor2   g1435(.a(G826), .b(n1274), .O(n1737));
  nor2   g1436(.a(n1269), .b(G164), .O(n1738));
  nor2   g1437(.a(G1691), .b(G194), .O(n1739));
  nor2   g1438(.a(n1739), .b(n1277), .O(n1740));
  inv1   g1439(.a(n1740), .O(n1741));
  nor2   g1440(.a(n1741), .b(n1738), .O(n1742));
  nor2   g1441(.a(n1742), .b(n1737), .O(n1743));
  inv1   g1442(.a(n1743), .O(n1744));
  nor2   g1443(.a(n1744), .b(n1736), .O(n1745));
  nor2   g1444(.a(n1745), .b(n1251), .O(G685));
  nor2   g1445(.a(G863), .b(n1271), .O(n1747));
  nor2   g1446(.a(G824), .b(n1274), .O(n1748));
  nor2   g1447(.a(n1269), .b(G161), .O(n1749));
  nor2   g1448(.a(G1691), .b(G191), .O(n1750));
  nor2   g1449(.a(n1750), .b(n1277), .O(n1751));
  inv1   g1450(.a(n1751), .O(n1752));
  nor2   g1451(.a(n1752), .b(n1749), .O(n1753));
  nor2   g1452(.a(n1753), .b(n1748), .O(n1754));
  inv1   g1453(.a(n1754), .O(n1755));
  nor2   g1454(.a(n1755), .b(n1747), .O(n1756));
  nor2   g1455(.a(n1756), .b(n1251), .O(G688));
  nor2   g1456(.a(n935), .b(G120), .O(n1758));
  nor2   g1457(.a(n813), .b(n787), .O(n1759));
  nor2   g1458(.a(n813), .b(n791), .O(n1760));
  nor2   g1459(.a(n796), .b(n788), .O(n1761));
  inv1   g1460(.a(n1761), .O(n1762));
  nor2   g1461(.a(n1762), .b(n1760), .O(n1763));
  nor2   g1462(.a(n1763), .b(n1759), .O(n1764));
  inv1   g1463(.a(n1764), .O(n1765));
  nor2   g1464(.a(n1032), .b(n805), .O(n1766));
  nor2   g1465(.a(n1031), .b(n804), .O(n1767));
  nor2   g1466(.a(n1767), .b(n1766), .O(n1768));
  inv1   g1467(.a(n1768), .O(n1769));
  nor2   g1468(.a(n1769), .b(n1765), .O(n1770));
  inv1   g1469(.a(G2174), .O(n1771));
  nor2   g1470(.a(n1768), .b(n1764), .O(n1772));
  nor2   g1471(.a(n1772), .b(n1771), .O(n1773));
  inv1   g1472(.a(n1773), .O(n1774));
  nor2   g1473(.a(n1774), .b(n1770), .O(n1775));
  inv1   g1474(.a(n813), .O(n1776));
  nor2   g1475(.a(n1776), .b(n804), .O(n1777));
  nor2   g1476(.a(n1777), .b(n814), .O(n1778));
  nor2   g1477(.a(n1032), .b(n789), .O(n1779));
  nor2   g1478(.a(n1779), .b(n791), .O(n1780));
  inv1   g1479(.a(n1780), .O(n1781));
  nor2   g1480(.a(n1781), .b(n1778), .O(n1782));
  inv1   g1481(.a(n1778), .O(n1783));
  nor2   g1482(.a(n1780), .b(n1783), .O(n1784));
  nor2   g1483(.a(n1784), .b(G2174), .O(n1785));
  inv1   g1484(.a(n1785), .O(n1786));
  nor2   g1485(.a(n1786), .b(n1782), .O(n1787));
  nor2   g1486(.a(n1787), .b(n1775), .O(n1788));
  nor2   g1487(.a(n817), .b(n1771), .O(n1789));
  nor2   g1488(.a(n1789), .b(n909), .O(n1790));
  inv1   g1489(.a(n1790), .O(n1791));
  nor2   g1490(.a(n915), .b(n739), .O(n1792));
  inv1   g1491(.a(n1792), .O(n1793));
  nor2   g1492(.a(n1793), .b(n743), .O(n1794));
  nor2   g1493(.a(n1792), .b(n1117), .O(n1795));
  nor2   g1494(.a(n1795), .b(n1794), .O(n1796));
  inv1   g1495(.a(n1796), .O(n1797));
  nor2   g1496(.a(n1797), .b(n1508), .O(n1798));
  nor2   g1497(.a(n1796), .b(n1509), .O(n1799));
  nor2   g1498(.a(n1799), .b(n1798), .O(n1800));
  nor2   g1499(.a(n1800), .b(n1791), .O(n1801));
  nor2   g1500(.a(n1797), .b(n765), .O(n1802));
  nor2   g1501(.a(n763), .b(n751), .O(n1803));
  nor2   g1502(.a(n1803), .b(n913), .O(n1804));
  inv1   g1503(.a(n1804), .O(n1805));
  nor2   g1504(.a(n983), .b(n766), .O(n1806));
  nor2   g1505(.a(n1806), .b(n1805), .O(n1807));
  inv1   g1506(.a(n1807), .O(n1808));
  nor2   g1507(.a(n1808), .b(n1802), .O(n1809));
  nor2   g1508(.a(n1804), .b(n1797), .O(n1810));
  nor2   g1509(.a(n1810), .b(n1809), .O(n1811));
  nor2   g1510(.a(n1811), .b(n1790), .O(n1812));
  nor2   g1511(.a(n1812), .b(n1801), .O(n1813));
  nor2   g1512(.a(n1813), .b(n969), .O(n1814));
  inv1   g1513(.a(n1813), .O(n1815));
  nor2   g1514(.a(n1815), .b(n968), .O(n1816));
  nor2   g1515(.a(n1816), .b(n1814), .O(n1817));
  nor2   g1516(.a(n1817), .b(n1788), .O(n1818));
  inv1   g1517(.a(n1788), .O(n1819));
  inv1   g1518(.a(n1817), .O(n1820));
  nor2   g1519(.a(n1820), .b(n1819), .O(n1821));
  nor2   g1520(.a(n1821), .b(n924), .O(n1822));
  inv1   g1521(.a(n1822), .O(n1823));
  nor2   g1522(.a(n1823), .b(n1818), .O(n1824));
  nor2   g1523(.a(n1516), .b(n1496), .O(n1825));
  nor2   g1524(.a(n1825), .b(n449), .O(n1826));
  inv1   g1525(.a(n1826), .O(n1827));
  nor2   g1526(.a(n398), .b(G248), .O(n1828));
  nor2   g1527(.a(G351), .b(G251), .O(n1829));
  nor2   g1528(.a(n1829), .b(n400), .O(n1830));
  inv1   g1529(.a(n1830), .O(n1831));
  nor2   g1530(.a(n1831), .b(n1828), .O(n1832));
  nor2   g1531(.a(n398), .b(n441), .O(n1833));
  nor2   g1532(.a(G351), .b(n443), .O(n1834));
  nor2   g1533(.a(n1834), .b(G534), .O(n1835));
  inv1   g1534(.a(n1835), .O(n1836));
  nor2   g1535(.a(n1836), .b(n1833), .O(n1837));
  nor2   g1536(.a(n1837), .b(n1832), .O(n1838));
  inv1   g1537(.a(n1838), .O(n1839));
  nor2   g1538(.a(n1839), .b(n463), .O(n1840));
  nor2   g1539(.a(n1838), .b(n1526), .O(n1841));
  nor2   g1540(.a(n1841), .b(n1840), .O(n1842));
  inv1   g1541(.a(n1842), .O(n1843));
  nor2   g1542(.a(G514), .b(G242), .O(n1844));
  nor2   g1543(.a(n475), .b(n428), .O(n1845));
  nor2   g1544(.a(n1845), .b(n1844), .O(n1846));
  nor2   g1545(.a(n1846), .b(n1843), .O(n1847));
  inv1   g1546(.a(n1846), .O(n1848));
  nor2   g1547(.a(n1848), .b(n1842), .O(n1849));
  nor2   g1548(.a(n1849), .b(n1847), .O(n1850));
  inv1   g1549(.a(n1850), .O(n1851));
  nor2   g1550(.a(n471), .b(n928), .O(n1852));
  nor2   g1551(.a(n1852), .b(n473), .O(n1853));
  nor2   g1552(.a(n411), .b(G248), .O(n1854));
  nor2   g1553(.a(G324), .b(G251), .O(n1855));
  nor2   g1554(.a(n1855), .b(n413), .O(n1856));
  inv1   g1555(.a(n1856), .O(n1857));
  nor2   g1556(.a(n1857), .b(n1854), .O(n1858));
  nor2   g1557(.a(n411), .b(n441), .O(n1859));
  nor2   g1558(.a(G324), .b(n443), .O(n1860));
  nor2   g1559(.a(n1860), .b(G503), .O(n1861));
  inv1   g1560(.a(n1861), .O(n1862));
  nor2   g1561(.a(n1862), .b(n1859), .O(n1863));
  nor2   g1562(.a(n1863), .b(n1858), .O(n1864));
  nor2   g1563(.a(n1864), .b(n1853), .O(n1865));
  inv1   g1564(.a(n1853), .O(n1866));
  inv1   g1565(.a(n1864), .O(n1867));
  nor2   g1566(.a(n1867), .b(n1866), .O(n1868));
  nor2   g1567(.a(n1868), .b(n1865), .O(n1869));
  inv1   g1568(.a(n1869), .O(n1870));
  nor2   g1569(.a(n383), .b(G248), .O(n1871));
  nor2   g1570(.a(G341), .b(G251), .O(n1872));
  nor2   g1571(.a(n1872), .b(n386), .O(n1873));
  inv1   g1572(.a(n1873), .O(n1874));
  nor2   g1573(.a(n1874), .b(n1871), .O(n1875));
  nor2   g1574(.a(n383), .b(n441), .O(n1876));
  nor2   g1575(.a(G341), .b(n443), .O(n1877));
  nor2   g1576(.a(n1877), .b(G523), .O(n1878));
  inv1   g1577(.a(n1878), .O(n1879));
  nor2   g1578(.a(n1879), .b(n1876), .O(n1880));
  nor2   g1579(.a(n1880), .b(n1875), .O(n1881));
  nor2   g1580(.a(n1881), .b(n1870), .O(n1882));
  inv1   g1581(.a(n1881), .O(n1883));
  nor2   g1582(.a(n1883), .b(n1869), .O(n1884));
  nor2   g1583(.a(n1884), .b(n1882), .O(n1885));
  inv1   g1584(.a(n1885), .O(n1886));
  nor2   g1585(.a(n1886), .b(n1851), .O(n1887));
  nor2   g1586(.a(n1885), .b(n1850), .O(n1888));
  nor2   g1587(.a(n1888), .b(n1887), .O(n1889));
  nor2   g1588(.a(n1889), .b(n1827), .O(n1890));
  inv1   g1589(.a(n1889), .O(n1891));
  nor2   g1590(.a(n1891), .b(n1826), .O(n1892));
  nor2   g1591(.a(n1892), .b(G4091), .O(n1893));
  inv1   g1592(.a(n1893), .O(n1894));
  nor2   g1593(.a(n1894), .b(n1890), .O(n1895));
  nor2   g1594(.a(n1895), .b(G4092), .O(n1896));
  inv1   g1595(.a(n1896), .O(n1897));
  nor2   g1596(.a(n1897), .b(n1824), .O(n1898));
  nor2   g1597(.a(n1898), .b(n1758), .O(G843));
  nor2   g1598(.a(n935), .b(G118), .O(n1900));
  inv1   g1599(.a(n896), .O(n1901));
  inv1   g1600(.a(G1497), .O(n1902));
  nor2   g1601(.a(n684), .b(n1902), .O(n1903));
  nor2   g1602(.a(n1903), .b(n1901), .O(n1904));
  inv1   g1603(.a(n1904), .O(n1905));
  inv1   g1604(.a(n712), .O(n1906));
  nor2   g1605(.a(n1906), .b(n692), .O(n1907));
  nor2   g1606(.a(n1907), .b(n713), .O(n1908));
  inv1   g1607(.a(n1908), .O(n1909));
  nor2   g1608(.a(n1193), .b(n689), .O(n1910));
  nor2   g1609(.a(n1910), .b(n899), .O(n1911));
  nor2   g1610(.a(n1911), .b(n723), .O(n1912));
  inv1   g1611(.a(n1911), .O(n1913));
  nor2   g1612(.a(n1913), .b(n722), .O(n1914));
  nor2   g1613(.a(n1914), .b(n1912), .O(n1915));
  inv1   g1614(.a(n1915), .O(n1916));
  nor2   g1615(.a(n1916), .b(n1909), .O(n1917));
  nor2   g1616(.a(n1915), .b(n1908), .O(n1918));
  nor2   g1617(.a(n1918), .b(n1917), .O(n1919));
  inv1   g1618(.a(n1919), .O(n1920));
  nor2   g1619(.a(n1920), .b(n1905), .O(n1921));
  nor2   g1620(.a(n728), .b(n722), .O(n1922));
  nor2   g1621(.a(n1922), .b(n730), .O(n1923));
  nor2   g1622(.a(n709), .b(n704), .O(n1924));
  inv1   g1623(.a(n1924), .O(n1925));
  nor2   g1624(.a(n1925), .b(n691), .O(n1926));
  nor2   g1625(.a(n1924), .b(n689), .O(n1927));
  nor2   g1626(.a(n1927), .b(n1926), .O(n1928));
  nor2   g1627(.a(n1928), .b(n1923), .O(n1929));
  inv1   g1628(.a(n1923), .O(n1930));
  inv1   g1629(.a(n1928), .O(n1931));
  nor2   g1630(.a(n1931), .b(n1930), .O(n1932));
  nor2   g1631(.a(n1932), .b(n1929), .O(n1933));
  inv1   g1632(.a(n1933), .O(n1934));
  nor2   g1633(.a(n1934), .b(n1904), .O(n1935));
  nor2   g1634(.a(n1935), .b(n1921), .O(n1936));
  inv1   g1635(.a(n894), .O(n1937));
  nor2   g1636(.a(n1937), .b(n681), .O(n1938));
  inv1   g1637(.a(n1938), .O(n1939));
  nor2   g1638(.a(n1939), .b(n645), .O(n1940));
  inv1   g1639(.a(n645), .O(n1941));
  nor2   g1640(.a(n1938), .b(n1941), .O(n1942));
  nor2   g1641(.a(n1942), .b(n1940), .O(n1943));
  inv1   g1642(.a(n1943), .O(n1944));
  nor2   g1643(.a(n891), .b(n667), .O(n1945));
  nor2   g1644(.a(n1945), .b(n640), .O(n1946));
  inv1   g1645(.a(n1945), .O(n1947));
  nor2   g1646(.a(n1947), .b(n639), .O(n1948));
  nor2   g1647(.a(n1948), .b(n1946), .O(n1949));
  inv1   g1648(.a(n1949), .O(n1950));
  nor2   g1649(.a(n1950), .b(n888), .O(n1951));
  nor2   g1650(.a(n1949), .b(n669), .O(n1952));
  nor2   g1651(.a(n1952), .b(n1951), .O(n1953));
  inv1   g1652(.a(n1953), .O(n1954));
  inv1   g1653(.a(n1218), .O(n1955));
  nor2   g1654(.a(n1955), .b(n657), .O(n1956));
  nor2   g1655(.a(n1218), .b(n658), .O(n1957));
  nor2   g1656(.a(n1957), .b(n1956), .O(n1958));
  nor2   g1657(.a(n1958), .b(n1954), .O(n1959));
  inv1   g1658(.a(n1958), .O(n1960));
  nor2   g1659(.a(n1960), .b(n1953), .O(n1961));
  nor2   g1660(.a(n1961), .b(n1959), .O(n1962));
  nor2   g1661(.a(n1962), .b(n1944), .O(n1963));
  inv1   g1662(.a(n1962), .O(n1964));
  nor2   g1663(.a(n1964), .b(n1943), .O(n1965));
  nor2   g1664(.a(n1965), .b(n1963), .O(n1966));
  nor2   g1665(.a(n1966), .b(n1902), .O(n1967));
  nor2   g1666(.a(n669), .b(n645), .O(n1968));
  nor2   g1667(.a(n1968), .b(n647), .O(n1969));
  inv1   g1668(.a(n1969), .O(n1970));
  inv1   g1669(.a(n892), .O(n1971));
  nor2   g1670(.a(n1971), .b(n674), .O(n1972));
  nor2   g1671(.a(n1972), .b(n893), .O(n1973));
  nor2   g1672(.a(n1973), .b(n640), .O(n1974));
  inv1   g1673(.a(n1973), .O(n1975));
  nor2   g1674(.a(n1975), .b(n639), .O(n1976));
  nor2   g1675(.a(n1976), .b(n1974), .O(n1977));
  inv1   g1676(.a(n1977), .O(n1978));
  nor2   g1677(.a(n1978), .b(n1970), .O(n1979));
  nor2   g1678(.a(n1977), .b(n1969), .O(n1980));
  nor2   g1679(.a(n1980), .b(n1979), .O(n1981));
  nor2   g1680(.a(n1219), .b(n658), .O(n1982));
  nor2   g1681(.a(n1220), .b(n657), .O(n1983));
  nor2   g1682(.a(n1983), .b(n1982), .O(n1984));
  inv1   g1683(.a(n1984), .O(n1985));
  nor2   g1684(.a(n1985), .b(n1981), .O(n1986));
  inv1   g1685(.a(n1981), .O(n1987));
  nor2   g1686(.a(n1984), .b(n1987), .O(n1988));
  nor2   g1687(.a(n1988), .b(n1986), .O(n1989));
  nor2   g1688(.a(n1989), .b(G1497), .O(n1990));
  nor2   g1689(.a(n1990), .b(n1967), .O(n1991));
  nor2   g1690(.a(n1991), .b(n678), .O(n1992));
  inv1   g1691(.a(n1991), .O(n1993));
  nor2   g1692(.a(n1993), .b(n677), .O(n1994));
  nor2   g1693(.a(n1994), .b(n1992), .O(n1995));
  nor2   g1694(.a(n1995), .b(n1936), .O(n1996));
  inv1   g1695(.a(n1936), .O(n1997));
  inv1   g1696(.a(n1995), .O(n1998));
  nor2   g1697(.a(n1998), .b(n1997), .O(n1999));
  nor2   g1698(.a(n1999), .b(n924), .O(n2000));
  inv1   g1699(.a(n2000), .O(n2001));
  nor2   g1700(.a(n2001), .b(n1996), .O(n2002));
  nor2   g1701(.a(n441), .b(n500), .O(n2003));
  nor2   g1702(.a(n443), .b(G210), .O(n2004));
  nor2   g1703(.a(n2004), .b(G457), .O(n2005));
  inv1   g1704(.a(n2005), .O(n2006));
  nor2   g1705(.a(n2006), .b(n2003), .O(n2007));
  nor2   g1706(.a(n508), .b(n428), .O(n2008));
  nor2   g1707(.a(n511), .b(n431), .O(n2009));
  nor2   g1708(.a(n2009), .b(n2008), .O(n2010));
  inv1   g1709(.a(n2010), .O(n2011));
  nor2   g1710(.a(n2011), .b(n2007), .O(n2012));
  inv1   g1711(.a(n2012), .O(n2013));
  nor2   g1712(.a(n441), .b(n608), .O(n2014));
  nor2   g1713(.a(n443), .b(G218), .O(n2015));
  nor2   g1714(.a(n2015), .b(G468), .O(n2016));
  inv1   g1715(.a(n2016), .O(n2017));
  nor2   g1716(.a(n2017), .b(n2014), .O(n2018));
  nor2   g1717(.a(n616), .b(n428), .O(n2019));
  nor2   g1718(.a(n619), .b(n431), .O(n2020));
  nor2   g1719(.a(n2020), .b(n2019), .O(n2021));
  inv1   g1720(.a(n2021), .O(n2022));
  nor2   g1721(.a(n2022), .b(n2018), .O(n2023));
  nor2   g1722(.a(n2023), .b(n2013), .O(n2024));
  inv1   g1723(.a(n2023), .O(n2025));
  nor2   g1724(.a(n2025), .b(n2012), .O(n2026));
  nor2   g1725(.a(n2026), .b(n2024), .O(n2027));
  nor2   g1726(.a(n516), .b(G248), .O(n2028));
  nor2   g1727(.a(G273), .b(G251), .O(n2029));
  nor2   g1728(.a(n2029), .b(n518), .O(n2030));
  inv1   g1729(.a(n2030), .O(n2031));
  nor2   g1730(.a(n2031), .b(n2028), .O(n2032));
  nor2   g1731(.a(n516), .b(n441), .O(n2033));
  nor2   g1732(.a(G273), .b(n443), .O(n2034));
  nor2   g1733(.a(n2034), .b(G411), .O(n2035));
  inv1   g1734(.a(n2035), .O(n2036));
  nor2   g1735(.a(n2036), .b(n2033), .O(n2037));
  nor2   g1736(.a(n2037), .b(n2032), .O(n2038));
  inv1   g1737(.a(n2038), .O(n2039));
  nor2   g1738(.a(n487), .b(G248), .O(n2040));
  nor2   g1739(.a(G265), .b(G251), .O(n2041));
  nor2   g1740(.a(n2041), .b(n489), .O(n2042));
  inv1   g1741(.a(n2042), .O(n2043));
  nor2   g1742(.a(n2043), .b(n2040), .O(n2044));
  nor2   g1743(.a(n487), .b(n441), .O(n2045));
  nor2   g1744(.a(G265), .b(n443), .O(n2046));
  nor2   g1745(.a(n2046), .b(G400), .O(n2047));
  inv1   g1746(.a(n2047), .O(n2048));
  nor2   g1747(.a(n2048), .b(n2045), .O(n2049));
  nor2   g1748(.a(n2049), .b(n2044), .O(n2050));
  inv1   g1749(.a(n2050), .O(n2051));
  nor2   g1750(.a(n441), .b(n577), .O(n2052));
  nor2   g1751(.a(n443), .b(G234), .O(n2053));
  nor2   g1752(.a(n2053), .b(G435), .O(n2054));
  inv1   g1753(.a(n2054), .O(n2055));
  nor2   g1754(.a(n2055), .b(n2052), .O(n2056));
  nor2   g1755(.a(n585), .b(n428), .O(n2057));
  nor2   g1756(.a(n588), .b(n431), .O(n2058));
  nor2   g1757(.a(n2058), .b(n2057), .O(n2059));
  inv1   g1758(.a(n2059), .O(n2060));
  nor2   g1759(.a(n2060), .b(n2056), .O(n2061));
  nor2   g1760(.a(n2061), .b(n2051), .O(n2062));
  inv1   g1761(.a(n2061), .O(n2063));
  nor2   g1762(.a(n2063), .b(n2050), .O(n2064));
  nor2   g1763(.a(n2064), .b(n2062), .O(n2065));
  nor2   g1764(.a(n2065), .b(n2039), .O(n2066));
  inv1   g1765(.a(n2065), .O(n2067));
  nor2   g1766(.a(n2067), .b(n2038), .O(n2068));
  nor2   g1767(.a(n2068), .b(n2066), .O(n2069));
  inv1   g1768(.a(n2069), .O(n2070));
  nor2   g1769(.a(n549), .b(G248), .O(n2071));
  nor2   g1770(.a(G281), .b(G251), .O(n2072));
  nor2   g1771(.a(n2072), .b(n551), .O(n2073));
  inv1   g1772(.a(n2073), .O(n2074));
  nor2   g1773(.a(n2074), .b(n2071), .O(n2075));
  nor2   g1774(.a(n549), .b(n441), .O(n2076));
  nor2   g1775(.a(G281), .b(n443), .O(n2077));
  nor2   g1776(.a(n2077), .b(G374), .O(n2078));
  inv1   g1777(.a(n2078), .O(n2079));
  nor2   g1778(.a(n2079), .b(n2076), .O(n2080));
  nor2   g1779(.a(n2080), .b(n2075), .O(n2081));
  inv1   g1780(.a(n2081), .O(n2082));
  nor2   g1781(.a(n564), .b(G248), .O(n2083));
  nor2   g1782(.a(G257), .b(G251), .O(n2084));
  nor2   g1783(.a(n2084), .b(n566), .O(n2085));
  inv1   g1784(.a(n2085), .O(n2086));
  nor2   g1785(.a(n2086), .b(n2083), .O(n2087));
  nor2   g1786(.a(n564), .b(n441), .O(n2088));
  nor2   g1787(.a(G257), .b(n443), .O(n2089));
  nor2   g1788(.a(n2089), .b(G389), .O(n2090));
  inv1   g1789(.a(n2090), .O(n2091));
  nor2   g1790(.a(n2091), .b(n2088), .O(n2092));
  nor2   g1791(.a(n2092), .b(n2087), .O(n2093));
  nor2   g1792(.a(n2093), .b(n1549), .O(n2094));
  inv1   g1793(.a(n2093), .O(n2095));
  nor2   g1794(.a(n2095), .b(n607), .O(n2096));
  nor2   g1795(.a(n2096), .b(n2094), .O(n2097));
  inv1   g1796(.a(n2097), .O(n2098));
  nor2   g1797(.a(n2098), .b(n2082), .O(n2099));
  nor2   g1798(.a(n2097), .b(n2081), .O(n2100));
  nor2   g1799(.a(n2100), .b(n2099), .O(n2101));
  inv1   g1800(.a(n2101), .O(n2102));
  nor2   g1801(.a(n441), .b(n533), .O(n2103));
  nor2   g1802(.a(n443), .b(G226), .O(n2104));
  nor2   g1803(.a(n2104), .b(G422), .O(n2105));
  inv1   g1804(.a(n2105), .O(n2106));
  nor2   g1805(.a(n2106), .b(n2103), .O(n2107));
  nor2   g1806(.a(n541), .b(n428), .O(n2108));
  nor2   g1807(.a(n544), .b(n431), .O(n2109));
  nor2   g1808(.a(n2109), .b(n2108), .O(n2110));
  inv1   g1809(.a(n2110), .O(n2111));
  nor2   g1810(.a(n2111), .b(n2107), .O(n2112));
  nor2   g1811(.a(n2112), .b(n2102), .O(n2113));
  inv1   g1812(.a(n2112), .O(n2114));
  nor2   g1813(.a(n2114), .b(n2101), .O(n2115));
  nor2   g1814(.a(n2115), .b(n2113), .O(n2116));
  inv1   g1815(.a(n2116), .O(n2117));
  nor2   g1816(.a(n2117), .b(n2070), .O(n2118));
  nor2   g1817(.a(n2116), .b(n2069), .O(n2119));
  nor2   g1818(.a(n2119), .b(n2118), .O(n2120));
  inv1   g1819(.a(n2120), .O(n2121));
  nor2   g1820(.a(n2121), .b(n2027), .O(n2122));
  inv1   g1821(.a(n2027), .O(n2123));
  nor2   g1822(.a(n2120), .b(n2123), .O(n2124));
  nor2   g1823(.a(n2124), .b(G4091), .O(n2125));
  inv1   g1824(.a(n2125), .O(n2126));
  nor2   g1825(.a(n2126), .b(n2122), .O(n2127));
  nor2   g1826(.a(n2127), .b(G4092), .O(n2128));
  inv1   g1827(.a(n2128), .O(n2129));
  nor2   g1828(.a(n2129), .b(n2002), .O(n2130));
  nor2   g1829(.a(n2130), .b(n1900), .O(G882));
  inv1   g1830(.a(G97), .O(n2132));
  nor2   g1831(.a(n933), .b(n2132), .O(n2133));
  nor2   g1832(.a(n2133), .b(n2130), .O(n2134));
  nor2   g1833(.a(n2134), .b(n989), .O(n2135));
  inv1   g1834(.a(G94), .O(n2136));
  nor2   g1835(.a(n933), .b(n2136), .O(n2137));
  nor2   g1836(.a(n2137), .b(n1898), .O(n2138));
  nor2   g1837(.a(n2138), .b(n992), .O(n2139));
  nor2   g1838(.a(n987), .b(G64), .O(n2140));
  nor2   g1839(.a(G4088), .b(G14), .O(n2141));
  nor2   g1840(.a(n2141), .b(n995), .O(n2142));
  inv1   g1841(.a(n2142), .O(n2143));
  nor2   g1842(.a(n2143), .b(n2140), .O(n2144));
  nor2   g1843(.a(n2144), .b(n2139), .O(n2145));
  inv1   g1844(.a(n2145), .O(n2146));
  nor2   g1845(.a(n2146), .b(n2135), .O(n2147));
  inv1   g1846(.a(n2147), .O(G767));
  nor2   g1847(.a(n2134), .b(n1046), .O(n2149));
  nor2   g1848(.a(n2138), .b(n1049), .O(n2150));
  nor2   g1849(.a(n1044), .b(G64), .O(n2151));
  nor2   g1850(.a(G4089), .b(G14), .O(n2152));
  nor2   g1851(.a(n2152), .b(n1052), .O(n2153));
  inv1   g1852(.a(n2153), .O(n2154));
  nor2   g1853(.a(n2154), .b(n2151), .O(n2155));
  nor2   g1854(.a(n2155), .b(n2150), .O(n2156));
  inv1   g1855(.a(n2156), .O(n2157));
  nor2   g1856(.a(n2157), .b(n2149), .O(n2158));
  inv1   g1857(.a(n2158), .O(G807));
  nor2   g1858(.a(n2134), .b(n1254), .O(n2160));
  nor2   g1859(.a(n2138), .b(n1257), .O(n2161));
  nor2   g1860(.a(n1252), .b(G179), .O(n2162));
  nor2   g1861(.a(G1689), .b(G176), .O(n2163));
  nor2   g1862(.a(n2163), .b(n1260), .O(n2164));
  inv1   g1863(.a(n2164), .O(n2165));
  nor2   g1864(.a(n2165), .b(n2162), .O(n2166));
  nor2   g1865(.a(n2166), .b(n2161), .O(n2167));
  inv1   g1866(.a(n2167), .O(n2168));
  nor2   g1867(.a(n2168), .b(n2160), .O(n2169));
  nor2   g1868(.a(n2169), .b(n1251), .O(n2170));
  inv1   g1869(.a(n2170), .O(G658));
  nor2   g1870(.a(n2134), .b(n1271), .O(n2172));
  nor2   g1871(.a(n2138), .b(n1274), .O(n2173));
  nor2   g1872(.a(n1269), .b(G179), .O(n2174));
  nor2   g1873(.a(G1691), .b(G176), .O(n2175));
  nor2   g1874(.a(n2175), .b(n1277), .O(n2176));
  inv1   g1875(.a(n2176), .O(n2177));
  nor2   g1876(.a(n2177), .b(n2174), .O(n2178));
  nor2   g1877(.a(n2178), .b(n2173), .O(n2179));
  inv1   g1878(.a(n2179), .O(n2180));
  nor2   g1879(.a(n2180), .b(n2172), .O(n2181));
  nor2   g1880(.a(n2181), .b(n1251), .O(n2182));
  inv1   g1881(.a(n2182), .O(G690));
  buffer g1882(.a(G141), .O(G144));
  buffer g1883(.a(G293), .O(G298));
  buffer g1884(.a(G3173), .O(G973));
  inv1   g1885(.a(G545), .O(G603));
  inv1   g1886(.a(G545), .O(G604));
  buffer g1887(.a(G137), .O(G926));
  buffer g1888(.a(G141), .O(G923));
  buffer g1889(.a(G1), .O(G921));
  buffer g1890(.a(G549), .O(G892));
  buffer g1891(.a(G299), .O(G887));
  inv1   g1892(.a(G549), .O(G606));
  buffer g1893(.a(G1), .O(G993));
  buffer g1894(.a(G1), .O(G978));
  buffer g1895(.a(G1), .O(G949));
  buffer g1896(.a(G1), .O(G939));
  buffer g1897(.a(G299), .O(G889));
  inv1   g1898(.a(n346), .O(G717));
  nor2   g1899(.a(n817), .b(n768), .O(G626));
  nor2   g1900(.a(n733), .b(n684), .O(G632));
  inv1   g1901(.a(n904), .O(G621));
  inv1   g1902(.a(n918), .O(G629));
endmodule


