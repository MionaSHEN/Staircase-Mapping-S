// Benchmark "c7552_blif" written by ABC on Sun Apr 14 20:30:20 2019

module c7552_blif  ( 
    G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47,
    G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65,
    G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83,
    G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110,
    G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133, G134,
    G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, G155, G156,
    G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, G167, G168,
    G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179, G180,
    G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G216,
    G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227, G228,
    G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239, G240,
    ING339 , G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492,
    G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247,
    G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737,
    G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427,
    G4432, G4437, G4526, G4528,
    G339, G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492,
    G490, G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552,
    G550, G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526,
    G524, G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446,
    G284, G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264,
    G270, G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416,
    G249, G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333,
    G336, G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471,
    G359, G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399  );
  input  G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41,
    G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63,
    G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81,
    G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106,
    G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130,
    G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154,
    G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166,
    G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190,
    G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202,
    G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214,
    G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226,
    G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238,
    G239, G240, ING339 , G1197, G1455, G1459, G1462, G1469, G1480, G1486,
    G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239,
    G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729,
    G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420,
    G4427, G4432, G4437, G4526, G4528;
  output G339, G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492,
    G490, G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552,
    G550, G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526,
    G524, G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446,
    G284, G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264,
    G270, G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416,
    G249, G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333,
    G336, G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471,
    G359, G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399;
  wire n317, n319, n320, n321, n322, n323, n324, n325, n326, n327, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n339, n340, n341, n342,
    n343, n344, n345, n346, n347, n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n359, n360, n362, n363, n364, n365, n366, n368, n369, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n869, n870, n871, n872, n873, n874, n875, n876, n877,
    n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
    n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
    n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
    n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
    n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
    n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
    n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
    n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
    n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
    n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
    n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
    n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
    n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
    n1358, n1359, n1360, n1361, n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1373, n1374, n1375, n1376, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386, n1388, n1389, n1390, n1392,
    n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
    n1403, n1404, n1405, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
    n1415, n1416, n1417, n1418, n1419, n1421, n1422, n1423, n1424, n1426,
    n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
    n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
    n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
    n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
    n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
    n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
    n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
    n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1766, n1767, n1768,
    n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
    n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
    n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
    n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
    n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
    n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
    n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1932, n1933, n1934, n1936, n1937, n1940, n1941, n1942,
    n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1951, n1952, n1953,
    n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1964, n1965,
    n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
    n1978, n1979, n1980, n1981, n1983, n1984, n1985, n1986, n1987, n1988,
    n1990, n1991, n1992, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2006, n2007, n2008, n2009, n2010, n2011,
    n2012, n2013, n2014, n2015, n2016, n2017, n2019, n2020, n2021, n2022,
    n2023, n2025, n2026, n2027, n2028, n2029, n2031, n2032, n2033, n2034,
    n2036, n2037, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
    n2048, n2049, n2050, n2051, n2052, n2053, n2055, n2056, n2057, n2058,
    n2059, n2060, n2061, n2062, n2063, n2064, n2066, n2067, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2080, n2081,
    n2082, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
    n2093, n2094, n2095, n2096, n2097, n2099, n2100, n2101, n2102, n2103,
    n2105, n2106, n2107, n2108, n2109, n2111, n2112, n2113, n2115, n2116,
    n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
    n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
    n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
    n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
    n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
    n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
    n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
    n2227, n2228, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
    n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
    n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
    n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
    n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
    n2308, n2309, n2310, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
    n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
    n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
    n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
    n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
    n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
    n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
    n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
    n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
    n2429, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
    n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
    n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
    n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
    n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
    n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
    n2540, n2541, n2542, n2543, n2544, n2545, n2546;
  inv1   g0000(.a(G15), .O(G279));
  nor2   g0001(.a(G57), .b(G5), .O(n317));
  inv1   g0002(.a(n317), .O(G402));
  inv1   g0003(.a(G228), .O(n319));
  inv1   g0004(.a(G240), .O(n320));
  nor2   g0005(.a(n320), .b(n319), .O(n321));
  inv1   g0006(.a(n321), .O(n322));
  inv1   g0007(.a(G150), .O(n323));
  inv1   g0008(.a(G184), .O(n324));
  nor2   g0009(.a(n324), .b(n323), .O(n325));
  inv1   g0010(.a(n325), .O(n326));
  nor2   g0011(.a(n326), .b(n322), .O(n327));
  inv1   g0012(.a(n327), .O(G404));
  inv1   g0013(.a(G218), .O(n329));
  inv1   g0014(.a(G230), .O(n330));
  nor2   g0015(.a(n330), .b(n329), .O(n331));
  inv1   g0016(.a(n331), .O(n332));
  inv1   g0017(.a(G152), .O(n333));
  inv1   g0018(.a(G210), .O(n334));
  nor2   g0019(.a(n334), .b(n333), .O(n335));
  inv1   g0020(.a(n335), .O(n336));
  nor2   g0021(.a(n336), .b(n332), .O(n337));
  inv1   g0022(.a(n337), .O(G406));
  inv1   g0023(.a(G185), .O(n339));
  inv1   g0024(.a(G186), .O(n340));
  nor2   g0025(.a(n340), .b(n339), .O(n341));
  inv1   g0026(.a(n341), .O(n342));
  inv1   g0027(.a(G182), .O(n343));
  inv1   g0028(.a(G183), .O(n344));
  nor2   g0029(.a(n344), .b(n343), .O(n345));
  inv1   g0030(.a(n345), .O(n346));
  nor2   g0031(.a(n346), .b(n342), .O(n347));
  inv1   g0032(.a(n347), .O(G408));
  inv1   g0033(.a(G188), .O(n349));
  inv1   g0034(.a(G199), .O(n350));
  nor2   g0035(.a(n350), .b(n349), .O(n351));
  inv1   g0036(.a(n351), .O(n352));
  inv1   g0037(.a(G162), .O(n353));
  inv1   g0038(.a(G172), .O(n354));
  nor2   g0039(.a(n354), .b(n353), .O(n355));
  inv1   g0040(.a(n355), .O(n356));
  nor2   g0041(.a(n356), .b(n352), .O(n357));
  inv1   g0042(.a(n357), .O(G410));
  inv1   g0043(.a(G1197), .O(n359));
  nor2   g0044(.a(n359), .b(G5), .O(n360));
  inv1   g0045(.a(n360), .O(G284));
  inv1   g0046(.a(G133), .O(n362));
  inv1   g0047(.a(G134), .O(n363));
  nor2   g0048(.a(n363), .b(n362), .O(n364));
  inv1   g0049(.a(n364), .O(n365));
  nor2   g0050(.a(n365), .b(G5), .O(n366));
  inv1   g0051(.a(n366), .O(G292));
  inv1   g0052(.a(G1), .O(n368));
  inv1   g0053(.a(G163), .O(n369));
  nor2   g0054(.a(n369), .b(n368), .O(G278));
  inv1   g0055(.a(G4526), .O(n371));
  inv1   g0056(.a(G41), .O(n372));
  nor2   g0057(.a(n372), .b(G18), .O(n373));
  inv1   g0058(.a(n373), .O(n374));
  nor2   g0059(.a(n374), .b(G3701), .O(n375));
  inv1   g0060(.a(G3701), .O(n376));
  nor2   g0061(.a(n376), .b(G18), .O(n377));
  inv1   g0062(.a(n377), .O(n378));
  nor2   g0063(.a(n378), .b(n373), .O(n379));
  nor2   g0064(.a(n379), .b(n375), .O(n380));
  inv1   g0065(.a(n380), .O(n381));
  nor2   g0066(.a(n381), .b(n371), .O(n382));
  nor2   g0067(.a(n380), .b(G4526), .O(n383));
  nor2   g0068(.a(n383), .b(n382), .O(G373));
  inv1   g0069(.a(G38), .O(n385));
  inv1   g0070(.a(G1492), .O(n386));
  inv1   g0071(.a(G4528), .O(n387));
  nor2   g0072(.a(n387), .b(n386), .O(n388));
  inv1   g0073(.a(n388), .O(n389));
  nor2   g0074(.a(n389), .b(n385), .O(n390));
  nor2   g0075(.a(n388), .b(G38), .O(n391));
  nor2   g0076(.a(n391), .b(n390), .O(n392));
  inv1   g0077(.a(G1496), .O(n393));
  nor2   g0078(.a(n387), .b(n393), .O(n394));
  nor2   g0079(.a(n394), .b(n385), .O(n395));
  nor2   g0080(.a(n387), .b(G38), .O(n396));
  inv1   g0081(.a(n396), .O(n397));
  nor2   g0082(.a(n397), .b(n393), .O(n398));
  nor2   g0083(.a(n398), .b(n395), .O(n399));
  inv1   g0084(.a(n399), .O(n400));
  nor2   g0085(.a(n400), .b(n392), .O(n401));
  inv1   g0086(.a(n401), .O(n402));
  inv1   g0087(.a(G9), .O(n403));
  inv1   g0088(.a(G12), .O(n404));
  nor2   g0089(.a(n404), .b(n403), .O(n405));
  inv1   g0090(.a(G18), .O(n406));
  nor2   g0091(.a(G213), .b(n406), .O(n407));
  nor2   g0092(.a(n407), .b(n405), .O(n408));
  inv1   g0093(.a(n408), .O(n409));
  nor2   g0094(.a(n409), .b(G1486), .O(n410));
  inv1   g0095(.a(G1486), .O(n411));
  nor2   g0096(.a(n408), .b(n411), .O(n412));
  nor2   g0097(.a(G214), .b(n406), .O(n413));
  nor2   g0098(.a(n413), .b(n405), .O(n414));
  inv1   g0099(.a(n414), .O(n415));
  nor2   g0100(.a(n415), .b(G1480), .O(n416));
  inv1   g0101(.a(n416), .O(n417));
  nor2   g0102(.a(n417), .b(n412), .O(n418));
  nor2   g0103(.a(n418), .b(n410), .O(n419));
  inv1   g0104(.a(n419), .O(n420));
  nor2   g0105(.a(n412), .b(n410), .O(n421));
  inv1   g0106(.a(n421), .O(n422));
  inv1   g0107(.a(G1480), .O(n423));
  nor2   g0108(.a(n414), .b(n423), .O(n424));
  nor2   g0109(.a(n424), .b(n416), .O(n425));
  inv1   g0110(.a(n425), .O(n426));
  nor2   g0111(.a(n426), .b(n422), .O(n427));
  inv1   g0112(.a(n427), .O(n428));
  nor2   g0113(.a(G209), .b(n406), .O(n429));
  nor2   g0114(.a(n429), .b(n405), .O(n430));
  inv1   g0115(.a(n430), .O(n431));
  nor2   g0116(.a(n431), .b(G1462), .O(n432));
  inv1   g0117(.a(n432), .O(n433));
  nor2   g0118(.a(G216), .b(n406), .O(n434));
  nor2   g0119(.a(n434), .b(n405), .O(n435));
  inv1   g0120(.a(n435), .O(n436));
  nor2   g0121(.a(n436), .b(G1469), .O(n437));
  inv1   g0122(.a(G1469), .O(n438));
  nor2   g0123(.a(n435), .b(n438), .O(n439));
  nor2   g0124(.a(n439), .b(n437), .O(n440));
  inv1   g0125(.a(n440), .O(n441));
  nor2   g0126(.a(n441), .b(n433), .O(n442));
  inv1   g0127(.a(n442), .O(n443));
  nor2   g0128(.a(G215), .b(n406), .O(n444));
  nor2   g0129(.a(n444), .b(n405), .O(n445));
  inv1   g0130(.a(n445), .O(n446));
  nor2   g0131(.a(n446), .b(G106), .O(n447));
  inv1   g0132(.a(G106), .O(n448));
  nor2   g0133(.a(n445), .b(n448), .O(n449));
  nor2   g0134(.a(n449), .b(n447), .O(n450));
  inv1   g0135(.a(n450), .O(n451));
  nor2   g0136(.a(n451), .b(n443), .O(n452));
  inv1   g0137(.a(n437), .O(n453));
  nor2   g0138(.a(n449), .b(n453), .O(n454));
  nor2   g0139(.a(n454), .b(n447), .O(n455));
  inv1   g0140(.a(n455), .O(n456));
  nor2   g0141(.a(n456), .b(n452), .O(n457));
  inv1   g0142(.a(n457), .O(n458));
  inv1   g0143(.a(G1462), .O(n459));
  nor2   g0144(.a(n430), .b(n459), .O(n460));
  nor2   g0145(.a(n460), .b(n432), .O(n461));
  inv1   g0146(.a(n461), .O(n462));
  nor2   g0147(.a(G154), .b(n406), .O(n463));
  nor2   g0148(.a(n463), .b(n405), .O(n464));
  inv1   g0149(.a(n464), .O(n465));
  nor2   g0150(.a(n465), .b(G2253), .O(n466));
  inv1   g0151(.a(G2253), .O(n467));
  nor2   g0152(.a(n464), .b(n467), .O(n468));
  nor2   g0153(.a(n468), .b(n466), .O(n469));
  inv1   g0154(.a(n469), .O(n470));
  inv1   g0155(.a(G2256), .O(n471));
  nor2   g0156(.a(G153), .b(n406), .O(n472));
  nor2   g0157(.a(n472), .b(n405), .O(n473));
  nor2   g0158(.a(n473), .b(n471), .O(n474));
  inv1   g0159(.a(n473), .O(n475));
  nor2   g0160(.a(n475), .b(G2256), .O(n476));
  nor2   g0161(.a(n476), .b(n474), .O(n477));
  inv1   g0162(.a(n477), .O(n478));
  nor2   g0163(.a(n478), .b(n470), .O(n479));
  inv1   g0164(.a(n479), .O(n480));
  nor2   g0165(.a(G156), .b(n406), .O(n481));
  nor2   g0166(.a(n481), .b(n405), .O(n482));
  inv1   g0167(.a(n482), .O(n483));
  nor2   g0168(.a(n483), .b(G2239), .O(n484));
  nor2   g0169(.a(G155), .b(n406), .O(n485));
  nor2   g0170(.a(n485), .b(n405), .O(n486));
  inv1   g0171(.a(n486), .O(n487));
  nor2   g0172(.a(n487), .b(G2247), .O(n488));
  inv1   g0173(.a(G2247), .O(n489));
  nor2   g0174(.a(n486), .b(n489), .O(n490));
  nor2   g0175(.a(n490), .b(n488), .O(n491));
  inv1   g0176(.a(n491), .O(n492));
  inv1   g0177(.a(G2239), .O(n493));
  nor2   g0178(.a(n482), .b(n493), .O(n494));
  nor2   g0179(.a(G157), .b(n406), .O(n495));
  nor2   g0180(.a(n495), .b(n405), .O(n496));
  inv1   g0181(.a(n496), .O(n497));
  nor2   g0182(.a(n497), .b(G2236), .O(n498));
  inv1   g0183(.a(G2236), .O(n499));
  nor2   g0184(.a(n496), .b(n499), .O(n500));
  nor2   g0185(.a(n500), .b(n498), .O(n501));
  inv1   g0186(.a(n501), .O(n502));
  inv1   g0187(.a(G135), .O(n503));
  nor2   g0188(.a(n503), .b(G18), .O(n504));
  inv1   g0189(.a(G158), .O(n505));
  nor2   g0190(.a(n505), .b(n406), .O(n506));
  nor2   g0191(.a(n506), .b(n504), .O(n507));
  nor2   g0192(.a(n507), .b(G2230), .O(n508));
  inv1   g0193(.a(G2230), .O(n509));
  inv1   g0194(.a(n507), .O(n510));
  nor2   g0195(.a(n510), .b(n509), .O(n511));
  nor2   g0196(.a(n511), .b(n508), .O(n512));
  inv1   g0197(.a(n512), .O(n513));
  nor2   g0198(.a(n513), .b(n502), .O(n514));
  inv1   g0199(.a(n514), .O(n515));
  inv1   g0200(.a(G2224), .O(n516));
  inv1   g0201(.a(G144), .O(n517));
  nor2   g0202(.a(n517), .b(G18), .O(n518));
  inv1   g0203(.a(G159), .O(n519));
  nor2   g0204(.a(n519), .b(n406), .O(n520));
  nor2   g0205(.a(n520), .b(n518), .O(n521));
  inv1   g0206(.a(n521), .O(n522));
  nor2   g0207(.a(n522), .b(n516), .O(n523));
  inv1   g0208(.a(G2218), .O(n524));
  inv1   g0209(.a(G138), .O(n525));
  nor2   g0210(.a(n525), .b(G18), .O(n526));
  inv1   g0211(.a(G160), .O(n527));
  nor2   g0212(.a(n527), .b(n406), .O(n528));
  nor2   g0213(.a(n528), .b(n526), .O(n529));
  inv1   g0214(.a(n529), .O(n530));
  nor2   g0215(.a(n530), .b(n524), .O(n531));
  inv1   g0216(.a(G147), .O(n532));
  nor2   g0217(.a(n532), .b(G18), .O(n533));
  inv1   g0218(.a(G151), .O(n534));
  nor2   g0219(.a(n534), .b(n406), .O(n535));
  nor2   g0220(.a(n535), .b(n533), .O(n536));
  nor2   g0221(.a(n536), .b(G2211), .O(n537));
  inv1   g0222(.a(n537), .O(n538));
  nor2   g0223(.a(n538), .b(n531), .O(n539));
  nor2   g0224(.a(n521), .b(G2224), .O(n540));
  nor2   g0225(.a(n529), .b(G2218), .O(n541));
  nor2   g0226(.a(n541), .b(n540), .O(n542));
  inv1   g0227(.a(n542), .O(n543));
  nor2   g0228(.a(n543), .b(n539), .O(n544));
  nor2   g0229(.a(n544), .b(n523), .O(n545));
  inv1   g0230(.a(n545), .O(n546));
  nor2   g0231(.a(n546), .b(n515), .O(n547));
  inv1   g0232(.a(n508), .O(n548));
  nor2   g0233(.a(n548), .b(n500), .O(n549));
  nor2   g0234(.a(n549), .b(n498), .O(n550));
  inv1   g0235(.a(n550), .O(n551));
  nor2   g0236(.a(n551), .b(n547), .O(n552));
  inv1   g0237(.a(n552), .O(n553));
  inv1   g0238(.a(G221), .O(n554));
  nor2   g0239(.a(n554), .b(n406), .O(n555));
  inv1   g0240(.a(G32), .O(n556));
  nor2   g0241(.a(n556), .b(G18), .O(n557));
  nor2   g0242(.a(n557), .b(n555), .O(n558));
  nor2   g0243(.a(n558), .b(G4427), .O(n559));
  inv1   g0244(.a(G4427), .O(n560));
  inv1   g0245(.a(n558), .O(n561));
  nor2   g0246(.a(n561), .b(n560), .O(n562));
  nor2   g0247(.a(n562), .b(n559), .O(n563));
  inv1   g0248(.a(n563), .O(n564));
  inv1   g0249(.a(G222), .O(n565));
  nor2   g0250(.a(n565), .b(n406), .O(n566));
  inv1   g0251(.a(G35), .O(n567));
  nor2   g0252(.a(n567), .b(G18), .O(n568));
  nor2   g0253(.a(n568), .b(n566), .O(n569));
  nor2   g0254(.a(n569), .b(G4420), .O(n570));
  inv1   g0255(.a(G4420), .O(n571));
  inv1   g0256(.a(n569), .O(n572));
  nor2   g0257(.a(n572), .b(n571), .O(n573));
  nor2   g0258(.a(n573), .b(n570), .O(n574));
  inv1   g0259(.a(n574), .O(n575));
  nor2   g0260(.a(n575), .b(n564), .O(n576));
  inv1   g0261(.a(n576), .O(n577));
  inv1   g0262(.a(G223), .O(n578));
  nor2   g0263(.a(n578), .b(n406), .O(n579));
  inv1   g0264(.a(G47), .O(n580));
  nor2   g0265(.a(n580), .b(G18), .O(n581));
  nor2   g0266(.a(n581), .b(n579), .O(n582));
  nor2   g0267(.a(n582), .b(G4415), .O(n583));
  inv1   g0268(.a(G4415), .O(n584));
  inv1   g0269(.a(n582), .O(n585));
  nor2   g0270(.a(n585), .b(n584), .O(n586));
  nor2   g0271(.a(n586), .b(n583), .O(n587));
  inv1   g0272(.a(n587), .O(n588));
  inv1   g0273(.a(G224), .O(n589));
  nor2   g0274(.a(n589), .b(n406), .O(n590));
  inv1   g0275(.a(G121), .O(n591));
  nor2   g0276(.a(n591), .b(G18), .O(n592));
  nor2   g0277(.a(n592), .b(n590), .O(n593));
  nor2   g0278(.a(n593), .b(G4410), .O(n594));
  inv1   g0279(.a(G4410), .O(n595));
  inv1   g0280(.a(n593), .O(n596));
  nor2   g0281(.a(n596), .b(n595), .O(n597));
  nor2   g0282(.a(n597), .b(n594), .O(n598));
  inv1   g0283(.a(n598), .O(n599));
  nor2   g0284(.a(n599), .b(n588), .O(n600));
  inv1   g0285(.a(n600), .O(n601));
  inv1   g0286(.a(G225), .O(n602));
  nor2   g0287(.a(n602), .b(n406), .O(n603));
  inv1   g0288(.a(G94), .O(n604));
  nor2   g0289(.a(n604), .b(G18), .O(n605));
  nor2   g0290(.a(n605), .b(n603), .O(n606));
  nor2   g0291(.a(n606), .b(G4405), .O(n607));
  inv1   g0292(.a(G226), .O(n608));
  nor2   g0293(.a(n608), .b(n406), .O(n609));
  inv1   g0294(.a(G97), .O(n610));
  nor2   g0295(.a(n610), .b(G18), .O(n611));
  nor2   g0296(.a(n611), .b(n609), .O(n612));
  nor2   g0297(.a(n612), .b(G4400), .O(n613));
  inv1   g0298(.a(n613), .O(n614));
  inv1   g0299(.a(G4405), .O(n615));
  inv1   g0300(.a(n606), .O(n616));
  nor2   g0301(.a(n616), .b(n615), .O(n617));
  nor2   g0302(.a(n617), .b(n614), .O(n618));
  nor2   g0303(.a(n618), .b(n607), .O(n619));
  inv1   g0304(.a(n619), .O(n620));
  inv1   g0305(.a(G217), .O(n621));
  nor2   g0306(.a(n621), .b(n406), .O(n622));
  inv1   g0307(.a(G118), .O(n623));
  nor2   g0308(.a(n623), .b(G18), .O(n624));
  nor2   g0309(.a(n624), .b(n622), .O(n625));
  nor2   g0310(.a(n625), .b(G4394), .O(n626));
  inv1   g0311(.a(n626), .O(n627));
  inv1   g0312(.a(G4400), .O(n628));
  inv1   g0313(.a(n612), .O(n629));
  nor2   g0314(.a(n629), .b(n628), .O(n630));
  nor2   g0315(.a(n630), .b(n613), .O(n631));
  inv1   g0316(.a(n631), .O(n632));
  nor2   g0317(.a(n632), .b(n627), .O(n633));
  inv1   g0318(.a(n633), .O(n634));
  nor2   g0319(.a(n617), .b(n607), .O(n635));
  inv1   g0320(.a(n635), .O(n636));
  nor2   g0321(.a(n636), .b(n634), .O(n637));
  nor2   g0322(.a(n637), .b(n620), .O(n638));
  nor2   g0323(.a(n638), .b(n601), .O(n639));
  nor2   g0324(.a(n594), .b(n583), .O(n640));
  nor2   g0325(.a(n640), .b(n586), .O(n641));
  nor2   g0326(.a(n641), .b(n639), .O(n642));
  inv1   g0327(.a(n642), .O(n643));
  inv1   g0328(.a(G4394), .O(n644));
  inv1   g0329(.a(n625), .O(n645));
  nor2   g0330(.a(n645), .b(n644), .O(n646));
  nor2   g0331(.a(n646), .b(n626), .O(n647));
  inv1   g0332(.a(n647), .O(n648));
  nor2   g0333(.a(n636), .b(n632), .O(n649));
  inv1   g0334(.a(n649), .O(n650));
  nor2   g0335(.a(n650), .b(n648), .O(n651));
  inv1   g0336(.a(n651), .O(n652));
  nor2   g0337(.a(n652), .b(n601), .O(n653));
  nor2   g0338(.a(n653), .b(n643), .O(n654));
  inv1   g0339(.a(G233), .O(n655));
  nor2   g0340(.a(n655), .b(n406), .O(n656));
  inv1   g0341(.a(G127), .O(n657));
  nor2   g0342(.a(n657), .b(G18), .O(n658));
  nor2   g0343(.a(n658), .b(n656), .O(n659));
  nor2   g0344(.a(n659), .b(G3737), .O(n660));
  inv1   g0345(.a(G3737), .O(n661));
  inv1   g0346(.a(n659), .O(n662));
  nor2   g0347(.a(n662), .b(n661), .O(n663));
  nor2   g0348(.a(n663), .b(n660), .O(n664));
  inv1   g0349(.a(n664), .O(n665));
  inv1   g0350(.a(G3729), .O(n666));
  inv1   g0351(.a(G234), .O(n667));
  nor2   g0352(.a(n667), .b(n406), .O(n668));
  inv1   g0353(.a(G130), .O(n669));
  nor2   g0354(.a(n669), .b(G18), .O(n670));
  nor2   g0355(.a(n670), .b(n668), .O(n671));
  inv1   g0356(.a(n671), .O(n672));
  nor2   g0357(.a(n672), .b(n666), .O(n673));
  inv1   g0358(.a(G235), .O(n674));
  nor2   g0359(.a(n674), .b(n406), .O(n675));
  inv1   g0360(.a(G103), .O(n676));
  nor2   g0361(.a(n676), .b(G18), .O(n677));
  nor2   g0362(.a(n677), .b(n675), .O(n678));
  nor2   g0363(.a(n678), .b(G3723), .O(n679));
  inv1   g0364(.a(G3723), .O(n680));
  inv1   g0365(.a(n678), .O(n681));
  nor2   g0366(.a(n681), .b(n680), .O(n682));
  nor2   g0367(.a(n682), .b(n679), .O(n683));
  inv1   g0368(.a(n683), .O(n684));
  inv1   g0369(.a(G236), .O(n685));
  nor2   g0370(.a(n685), .b(n406), .O(n686));
  inv1   g0371(.a(G23), .O(n687));
  nor2   g0372(.a(n687), .b(G18), .O(n688));
  nor2   g0373(.a(n688), .b(n686), .O(n689));
  nor2   g0374(.a(n689), .b(G3717), .O(n690));
  inv1   g0375(.a(G3717), .O(n691));
  inv1   g0376(.a(n689), .O(n692));
  nor2   g0377(.a(n692), .b(n691), .O(n693));
  nor2   g0378(.a(n693), .b(n690), .O(n694));
  inv1   g0379(.a(n694), .O(n695));
  nor2   g0380(.a(n695), .b(n684), .O(n696));
  inv1   g0381(.a(n696), .O(n697));
  inv1   g0382(.a(G3711), .O(n698));
  inv1   g0383(.a(G237), .O(n699));
  nor2   g0384(.a(n699), .b(n406), .O(n700));
  inv1   g0385(.a(G26), .O(n701));
  nor2   g0386(.a(n701), .b(G18), .O(n702));
  nor2   g0387(.a(n702), .b(n700), .O(n703));
  inv1   g0388(.a(n703), .O(n704));
  nor2   g0389(.a(n704), .b(n698), .O(n705));
  nor2   g0390(.a(n703), .b(G3711), .O(n706));
  inv1   g0391(.a(G238), .O(n707));
  nor2   g0392(.a(n707), .b(n406), .O(n708));
  inv1   g0393(.a(G29), .O(n709));
  nor2   g0394(.a(n709), .b(G18), .O(n710));
  nor2   g0395(.a(n710), .b(n708), .O(n711));
  nor2   g0396(.a(n711), .b(G3705), .O(n712));
  nor2   g0397(.a(n712), .b(n706), .O(n713));
  nor2   g0398(.a(n713), .b(n705), .O(n714));
  inv1   g0399(.a(n714), .O(n715));
  nor2   g0400(.a(n715), .b(n697), .O(n716));
  inv1   g0401(.a(n375), .O(n717));
  nor2   g0402(.a(n706), .b(n705), .O(n718));
  inv1   g0403(.a(n718), .O(n719));
  inv1   g0404(.a(G3705), .O(n720));
  inv1   g0405(.a(n711), .O(n721));
  nor2   g0406(.a(n721), .b(n720), .O(n722));
  nor2   g0407(.a(n722), .b(n712), .O(n723));
  inv1   g0408(.a(n723), .O(n724));
  nor2   g0409(.a(n724), .b(n719), .O(n725));
  inv1   g0410(.a(n725), .O(n726));
  nor2   g0411(.a(n726), .b(n717), .O(n727));
  inv1   g0412(.a(n727), .O(n728));
  nor2   g0413(.a(n728), .b(n693), .O(n729));
  nor2   g0414(.a(n729), .b(n690), .O(n730));
  inv1   g0415(.a(n730), .O(n731));
  nor2   g0416(.a(n731), .b(n679), .O(n732));
  nor2   g0417(.a(n732), .b(n682), .O(n733));
  nor2   g0418(.a(n733), .b(n716), .O(n734));
  inv1   g0419(.a(n734), .O(n735));
  nor2   g0420(.a(n726), .b(n381), .O(n736));
  inv1   g0421(.a(n736), .O(n737));
  nor2   g0422(.a(n737), .b(n697), .O(n738));
  inv1   g0423(.a(n738), .O(n739));
  nor2   g0424(.a(n739), .b(n371), .O(n740));
  nor2   g0425(.a(n740), .b(n735), .O(n741));
  nor2   g0426(.a(n741), .b(n673), .O(n742));
  inv1   g0427(.a(n742), .O(n743));
  nor2   g0428(.a(n743), .b(n665), .O(n744));
  inv1   g0429(.a(n744), .O(n745));
  nor2   g0430(.a(n671), .b(G3729), .O(n746));
  inv1   g0431(.a(G231), .O(n747));
  nor2   g0432(.a(n747), .b(n406), .O(n748));
  inv1   g0433(.a(G100), .O(n749));
  nor2   g0434(.a(n749), .b(G18), .O(n750));
  nor2   g0435(.a(n750), .b(n748), .O(n751));
  nor2   g0436(.a(n751), .b(G3749), .O(n752));
  inv1   g0437(.a(G3749), .O(n753));
  inv1   g0438(.a(n751), .O(n754));
  nor2   g0439(.a(n754), .b(n753), .O(n755));
  nor2   g0440(.a(n755), .b(n752), .O(n756));
  inv1   g0441(.a(n756), .O(n757));
  inv1   g0442(.a(G232), .O(n758));
  nor2   g0443(.a(n758), .b(n406), .O(n759));
  inv1   g0444(.a(G124), .O(n760));
  nor2   g0445(.a(n760), .b(G18), .O(n761));
  nor2   g0446(.a(n761), .b(n759), .O(n762));
  nor2   g0447(.a(n762), .b(G3743), .O(n763));
  inv1   g0448(.a(G3743), .O(n764));
  inv1   g0449(.a(n762), .O(n765));
  nor2   g0450(.a(n765), .b(n764), .O(n766));
  nor2   g0451(.a(n766), .b(n763), .O(n767));
  inv1   g0452(.a(n767), .O(n768));
  nor2   g0453(.a(n768), .b(n757), .O(n769));
  inv1   g0454(.a(n769), .O(n770));
  nor2   g0455(.a(n770), .b(n746), .O(n771));
  inv1   g0456(.a(n771), .O(n772));
  nor2   g0457(.a(n772), .b(n745), .O(n773));
  inv1   g0458(.a(n746), .O(n774));
  nor2   g0459(.a(n774), .b(n665), .O(n775));
  nor2   g0460(.a(n775), .b(n660), .O(n776));
  nor2   g0461(.a(n776), .b(n766), .O(n777));
  nor2   g0462(.a(n777), .b(n763), .O(n778));
  nor2   g0463(.a(n778), .b(n755), .O(n779));
  nor2   g0464(.a(n779), .b(n752), .O(n780));
  inv1   g0465(.a(n780), .O(n781));
  nor2   g0466(.a(n781), .b(n773), .O(n782));
  inv1   g0467(.a(n782), .O(n783));
  nor2   g0468(.a(n783), .b(n643), .O(n784));
  nor2   g0469(.a(n784), .b(n654), .O(n785));
  inv1   g0470(.a(n785), .O(n786));
  nor2   g0471(.a(n786), .b(n577), .O(n787));
  inv1   g0472(.a(n787), .O(n788));
  inv1   g0473(.a(G220), .O(n789));
  nor2   g0474(.a(n789), .b(n406), .O(n790));
  inv1   g0475(.a(G50), .O(n791));
  nor2   g0476(.a(n791), .b(G18), .O(n792));
  nor2   g0477(.a(n792), .b(n790), .O(n793));
  nor2   g0478(.a(n793), .b(G4432), .O(n794));
  inv1   g0479(.a(G4432), .O(n795));
  inv1   g0480(.a(n793), .O(n796));
  nor2   g0481(.a(n796), .b(n795), .O(n797));
  nor2   g0482(.a(n797), .b(n794), .O(n798));
  inv1   g0483(.a(n798), .O(n799));
  inv1   g0484(.a(G4437), .O(n800));
  inv1   g0485(.a(G219), .O(n801));
  nor2   g0486(.a(n801), .b(n406), .O(n802));
  inv1   g0487(.a(G66), .O(n803));
  nor2   g0488(.a(n803), .b(G18), .O(n804));
  nor2   g0489(.a(n804), .b(n802), .O(n805));
  inv1   g0490(.a(n805), .O(n806));
  nor2   g0491(.a(n806), .b(n800), .O(n807));
  nor2   g0492(.a(n805), .b(G4437), .O(n808));
  nor2   g0493(.a(n808), .b(n807), .O(n809));
  inv1   g0494(.a(n809), .O(n810));
  nor2   g0495(.a(n810), .b(n799), .O(n811));
  inv1   g0496(.a(n811), .O(n812));
  nor2   g0497(.a(n812), .b(n788), .O(n813));
  nor2   g0498(.a(n570), .b(n559), .O(n814));
  nor2   g0499(.a(n814), .b(n562), .O(n815));
  nor2   g0500(.a(n815), .b(n794), .O(n816));
  nor2   g0501(.a(n816), .b(n797), .O(n817));
  nor2   g0502(.a(n817), .b(n808), .O(n818));
  nor2   g0503(.a(n818), .b(n807), .O(n819));
  nor2   g0504(.a(n819), .b(n813), .O(n820));
  nor2   g0505(.a(n540), .b(n523), .O(n821));
  inv1   g0506(.a(n821), .O(n822));
  nor2   g0507(.a(n541), .b(n531), .O(n823));
  inv1   g0508(.a(n823), .O(n824));
  inv1   g0509(.a(G2211), .O(n825));
  inv1   g0510(.a(n536), .O(n826));
  nor2   g0511(.a(n826), .b(n825), .O(n827));
  nor2   g0512(.a(n827), .b(n537), .O(n828));
  inv1   g0513(.a(n828), .O(n829));
  nor2   g0514(.a(n829), .b(n824), .O(n830));
  inv1   g0515(.a(n830), .O(n831));
  nor2   g0516(.a(n831), .b(n822), .O(n832));
  inv1   g0517(.a(n832), .O(n833));
  nor2   g0518(.a(n833), .b(n515), .O(n834));
  inv1   g0519(.a(n834), .O(n835));
  nor2   g0520(.a(n835), .b(n820), .O(n836));
  nor2   g0521(.a(n836), .b(n553), .O(n837));
  nor2   g0522(.a(n837), .b(n494), .O(n838));
  inv1   g0523(.a(n838), .O(n839));
  nor2   g0524(.a(n839), .b(n492), .O(n840));
  inv1   g0525(.a(n840), .O(n841));
  nor2   g0526(.a(n841), .b(n484), .O(n842));
  inv1   g0527(.a(n842), .O(n843));
  nor2   g0528(.a(n843), .b(n480), .O(n844));
  inv1   g0529(.a(n484), .O(n845));
  nor2   g0530(.a(n492), .b(n845), .O(n846));
  nor2   g0531(.a(n846), .b(n488), .O(n847));
  inv1   g0532(.a(n847), .O(n848));
  nor2   g0533(.a(n848), .b(n466), .O(n849));
  nor2   g0534(.a(n849), .b(n468), .O(n850));
  nor2   g0535(.a(n850), .b(n476), .O(n851));
  nor2   g0536(.a(n851), .b(n474), .O(n852));
  nor2   g0537(.a(n852), .b(n844), .O(n853));
  nor2   g0538(.a(n853), .b(n462), .O(n854));
  inv1   g0539(.a(n854), .O(n855));
  nor2   g0540(.a(n855), .b(n441), .O(n856));
  inv1   g0541(.a(n856), .O(n857));
  nor2   g0542(.a(n857), .b(n451), .O(n858));
  nor2   g0543(.a(n858), .b(n458), .O(n859));
  nor2   g0544(.a(n859), .b(n428), .O(n860));
  nor2   g0545(.a(n860), .b(n420), .O(n861));
  nor2   g0546(.a(n861), .b(n402), .O(n862));
  nor2   g0547(.a(n388), .b(n385), .O(n863));
  nor2   g0548(.a(G1496), .b(n385), .O(n864));
  nor2   g0549(.a(n864), .b(n863), .O(n865));
  inv1   g0550(.a(n865), .O(n866));
  nor2   g0551(.a(n866), .b(n862), .O(n867));
  inv1   g0552(.a(n867), .O(G246));
  inv1   g0553(.a(G1455), .O(n869));
  inv1   g0554(.a(G2204), .O(n870));
  nor2   g0555(.a(n870), .b(n869), .O(n871));
  nor2   g0556(.a(n871), .b(n397), .O(n872));
  nor2   g0557(.a(G166), .b(n406), .O(n873));
  nor2   g0558(.a(n873), .b(n405), .O(n874));
  nor2   g0559(.a(n411), .b(n406), .O(n875));
  nor2   g0560(.a(G88), .b(G18), .O(n876));
  nor2   g0561(.a(n876), .b(n875), .O(n877));
  nor2   g0562(.a(n877), .b(n874), .O(n878));
  nor2   g0563(.a(G167), .b(n406), .O(n879));
  nor2   g0564(.a(n879), .b(n405), .O(n880));
  inv1   g0565(.a(n880), .O(n881));
  nor2   g0566(.a(n423), .b(n406), .O(n882));
  nor2   g0567(.a(G112), .b(G18), .O(n883));
  nor2   g0568(.a(n883), .b(n882), .O(n884));
  inv1   g0569(.a(n884), .O(n885));
  nor2   g0570(.a(n885), .b(n881), .O(n886));
  nor2   g0571(.a(G168), .b(n406), .O(n887));
  nor2   g0572(.a(n887), .b(n405), .O(n888));
  inv1   g0573(.a(n888), .O(n889));
  nor2   g0574(.a(n448), .b(n406), .O(n890));
  nor2   g0575(.a(G87), .b(G18), .O(n891));
  nor2   g0576(.a(n891), .b(n890), .O(n892));
  inv1   g0577(.a(n892), .O(n893));
  nor2   g0578(.a(n893), .b(n889), .O(n894));
  nor2   g0579(.a(n892), .b(n888), .O(n895));
  nor2   g0580(.a(n895), .b(n894), .O(n896));
  inv1   g0581(.a(n896), .O(n897));
  nor2   g0582(.a(G169), .b(n406), .O(n898));
  nor2   g0583(.a(n898), .b(n405), .O(n899));
  inv1   g0584(.a(n899), .O(n900));
  nor2   g0585(.a(n438), .b(n406), .O(n901));
  nor2   g0586(.a(G111), .b(G18), .O(n902));
  nor2   g0587(.a(n902), .b(n901), .O(n903));
  inv1   g0588(.a(n903), .O(n904));
  nor2   g0589(.a(n904), .b(n900), .O(n905));
  nor2   g0590(.a(n903), .b(n899), .O(n906));
  nor2   g0591(.a(n906), .b(n905), .O(n907));
  inv1   g0592(.a(n907), .O(n908));
  nor2   g0593(.a(n908), .b(n897), .O(n909));
  inv1   g0594(.a(n909), .O(n910));
  nor2   g0595(.a(n884), .b(n880), .O(n911));
  nor2   g0596(.a(n459), .b(n406), .O(n912));
  nor2   g0597(.a(G113), .b(G18), .O(n913));
  nor2   g0598(.a(n913), .b(n912), .O(n914));
  inv1   g0599(.a(n914), .O(n915));
  nor2   g0600(.a(n915), .b(n405), .O(n916));
  inv1   g0601(.a(n916), .O(n917));
  nor2   g0602(.a(n917), .b(n911), .O(n918));
  inv1   g0603(.a(n918), .O(n919));
  nor2   g0604(.a(n919), .b(n910), .O(n920));
  nor2   g0605(.a(n920), .b(n886), .O(n921));
  nor2   g0606(.a(n921), .b(n878), .O(n922));
  inv1   g0607(.a(G192), .O(n923));
  nor2   g0608(.a(n923), .b(n406), .O(n924));
  nor2   g0609(.a(n924), .b(n568), .O(n925));
  nor2   g0610(.a(n571), .b(n406), .O(n926));
  nor2   g0611(.a(G79), .b(G18), .O(n927));
  nor2   g0612(.a(n927), .b(n926), .O(n928));
  inv1   g0613(.a(n928), .O(n929));
  nor2   g0614(.a(n929), .b(n925), .O(n930));
  inv1   g0615(.a(G191), .O(n931));
  nor2   g0616(.a(n931), .b(n406), .O(n932));
  nor2   g0617(.a(n932), .b(n557), .O(n933));
  nor2   g0618(.a(n560), .b(n406), .O(n934));
  nor2   g0619(.a(G60), .b(G18), .O(n935));
  nor2   g0620(.a(n935), .b(n934), .O(n936));
  inv1   g0621(.a(n936), .O(n937));
  nor2   g0622(.a(n937), .b(n933), .O(n938));
  nor2   g0623(.a(n938), .b(n930), .O(n939));
  inv1   g0624(.a(G190), .O(n940));
  nor2   g0625(.a(n940), .b(n406), .O(n941));
  nor2   g0626(.a(n941), .b(n792), .O(n942));
  nor2   g0627(.a(n795), .b(n406), .O(n943));
  nor2   g0628(.a(G61), .b(G18), .O(n944));
  nor2   g0629(.a(n944), .b(n943), .O(n945));
  inv1   g0630(.a(n945), .O(n946));
  nor2   g0631(.a(n946), .b(n942), .O(n947));
  inv1   g0632(.a(n942), .O(n948));
  nor2   g0633(.a(n945), .b(n948), .O(n949));
  nor2   g0634(.a(n949), .b(n947), .O(n950));
  inv1   g0635(.a(n950), .O(n951));
  inv1   g0636(.a(n933), .O(n952));
  nor2   g0637(.a(n936), .b(n952), .O(n953));
  inv1   g0638(.a(G189), .O(n954));
  nor2   g0639(.a(n954), .b(n406), .O(n955));
  nor2   g0640(.a(n955), .b(n804), .O(n956));
  inv1   g0641(.a(n956), .O(n957));
  nor2   g0642(.a(n800), .b(n406), .O(n958));
  nor2   g0643(.a(G62), .b(G18), .O(n959));
  nor2   g0644(.a(n959), .b(n958), .O(n960));
  nor2   g0645(.a(n960), .b(n957), .O(n961));
  inv1   g0646(.a(n960), .O(n962));
  nor2   g0647(.a(n962), .b(n956), .O(n963));
  nor2   g0648(.a(n963), .b(n961), .O(n964));
  inv1   g0649(.a(n964), .O(n965));
  nor2   g0650(.a(n965), .b(n953), .O(n966));
  inv1   g0651(.a(n966), .O(n967));
  nor2   g0652(.a(n967), .b(n951), .O(n968));
  inv1   g0653(.a(n968), .O(n969));
  nor2   g0654(.a(n969), .b(n939), .O(n970));
  inv1   g0655(.a(n939), .O(n971));
  inv1   g0656(.a(n925), .O(n972));
  nor2   g0657(.a(n928), .b(n972), .O(n973));
  nor2   g0658(.a(n973), .b(n971), .O(n974));
  inv1   g0659(.a(n974), .O(n975));
  nor2   g0660(.a(n975), .b(n969), .O(n976));
  inv1   g0661(.a(n976), .O(n977));
  inv1   g0662(.a(G200), .O(n978));
  nor2   g0663(.a(n978), .b(n406), .O(n979));
  nor2   g0664(.a(n979), .b(n750), .O(n980));
  nor2   g0665(.a(n753), .b(n406), .O(n981));
  nor2   g0666(.a(G56), .b(G18), .O(n982));
  nor2   g0667(.a(n982), .b(n981), .O(n983));
  inv1   g0668(.a(n983), .O(n984));
  nor2   g0669(.a(n984), .b(n980), .O(n985));
  inv1   g0670(.a(G202), .O(n986));
  nor2   g0671(.a(n986), .b(n406), .O(n987));
  nor2   g0672(.a(n987), .b(n658), .O(n988));
  inv1   g0673(.a(n988), .O(n989));
  nor2   g0674(.a(n661), .b(n406), .O(n990));
  nor2   g0675(.a(G54), .b(G18), .O(n991));
  nor2   g0676(.a(n991), .b(n990), .O(n992));
  nor2   g0677(.a(n992), .b(n989), .O(n993));
  inv1   g0678(.a(n980), .O(n994));
  nor2   g0679(.a(n983), .b(n994), .O(n995));
  nor2   g0680(.a(n995), .b(n985), .O(n996));
  inv1   g0681(.a(n996), .O(n997));
  nor2   g0682(.a(n997), .b(n993), .O(n998));
  inv1   g0683(.a(n998), .O(n999));
  inv1   g0684(.a(n992), .O(n1000));
  nor2   g0685(.a(n1000), .b(n988), .O(n1001));
  inv1   g0686(.a(G203), .O(n1002));
  nor2   g0687(.a(n1002), .b(n406), .O(n1003));
  nor2   g0688(.a(n1003), .b(n670), .O(n1004));
  nor2   g0689(.a(n666), .b(n406), .O(n1005));
  nor2   g0690(.a(G53), .b(G18), .O(n1006));
  nor2   g0691(.a(n1006), .b(n1005), .O(n1007));
  inv1   g0692(.a(n1007), .O(n1008));
  nor2   g0693(.a(n1008), .b(n1004), .O(n1009));
  inv1   g0694(.a(G204), .O(n1010));
  nor2   g0695(.a(n1010), .b(n406), .O(n1011));
  nor2   g0696(.a(n1011), .b(n677), .O(n1012));
  inv1   g0697(.a(n1012), .O(n1013));
  nor2   g0698(.a(n680), .b(n406), .O(n1014));
  nor2   g0699(.a(G73), .b(G18), .O(n1015));
  nor2   g0700(.a(n1015), .b(n1014), .O(n1016));
  nor2   g0701(.a(n1016), .b(n1013), .O(n1017));
  nor2   g0702(.a(G89), .b(G70), .O(n1018));
  inv1   g0703(.a(G207), .O(n1019));
  nor2   g0704(.a(n1019), .b(n406), .O(n1020));
  nor2   g0705(.a(n1020), .b(n710), .O(n1021));
  inv1   g0706(.a(n1021), .O(n1022));
  nor2   g0707(.a(n720), .b(n406), .O(n1023));
  nor2   g0708(.a(G74), .b(G18), .O(n1024));
  nor2   g0709(.a(n1024), .b(n1023), .O(n1025));
  nor2   g0710(.a(n1025), .b(n1022), .O(n1026));
  inv1   g0711(.a(G89), .O(n1027));
  nor2   g0712(.a(G70), .b(G18), .O(n1028));
  nor2   g0713(.a(n1028), .b(n1027), .O(n1029));
  nor2   g0714(.a(n1029), .b(n373), .O(n1030));
  nor2   g0715(.a(n1030), .b(n1026), .O(n1031));
  inv1   g0716(.a(n1031), .O(n1032));
  nor2   g0717(.a(n1032), .b(n1018), .O(n1033));
  inv1   g0718(.a(G206), .O(n1034));
  nor2   g0719(.a(n1034), .b(n406), .O(n1035));
  nor2   g0720(.a(n1035), .b(n702), .O(n1036));
  nor2   g0721(.a(n698), .b(n406), .O(n1037));
  nor2   g0722(.a(G76), .b(G18), .O(n1038));
  nor2   g0723(.a(n1038), .b(n1037), .O(n1039));
  inv1   g0724(.a(n1039), .O(n1040));
  nor2   g0725(.a(n1040), .b(n1036), .O(n1041));
  inv1   g0726(.a(n1025), .O(n1042));
  nor2   g0727(.a(n1042), .b(n1021), .O(n1043));
  nor2   g0728(.a(n1043), .b(n1041), .O(n1044));
  inv1   g0729(.a(n1044), .O(n1045));
  nor2   g0730(.a(n1045), .b(n1033), .O(n1046));
  inv1   g0731(.a(G205), .O(n1047));
  nor2   g0732(.a(n1047), .b(n406), .O(n1048));
  nor2   g0733(.a(n1048), .b(n688), .O(n1049));
  inv1   g0734(.a(n1049), .O(n1050));
  nor2   g0735(.a(n691), .b(n406), .O(n1051));
  nor2   g0736(.a(G75), .b(G18), .O(n1052));
  nor2   g0737(.a(n1052), .b(n1051), .O(n1053));
  nor2   g0738(.a(n1053), .b(n1050), .O(n1054));
  inv1   g0739(.a(n1036), .O(n1055));
  nor2   g0740(.a(n1039), .b(n1055), .O(n1056));
  nor2   g0741(.a(n1056), .b(n1054), .O(n1057));
  inv1   g0742(.a(n1057), .O(n1058));
  nor2   g0743(.a(n1058), .b(n1046), .O(n1059));
  inv1   g0744(.a(n1016), .O(n1060));
  nor2   g0745(.a(n1060), .b(n1012), .O(n1061));
  inv1   g0746(.a(n1053), .O(n1062));
  nor2   g0747(.a(n1062), .b(n1049), .O(n1063));
  nor2   g0748(.a(n1063), .b(n1061), .O(n1064));
  inv1   g0749(.a(n1064), .O(n1065));
  nor2   g0750(.a(n1065), .b(n1059), .O(n1066));
  inv1   g0751(.a(n1004), .O(n1067));
  nor2   g0752(.a(n1007), .b(n1067), .O(n1068));
  nor2   g0753(.a(n1068), .b(n1066), .O(n1069));
  inv1   g0754(.a(n1069), .O(n1070));
  nor2   g0755(.a(n1070), .b(n1017), .O(n1071));
  nor2   g0756(.a(n1071), .b(n1009), .O(n1072));
  inv1   g0757(.a(n1072), .O(n1073));
  nor2   g0758(.a(n1073), .b(n1001), .O(n1074));
  inv1   g0759(.a(G201), .O(n1075));
  nor2   g0760(.a(n1075), .b(n406), .O(n1076));
  nor2   g0761(.a(n1076), .b(n761), .O(n1077));
  nor2   g0762(.a(n764), .b(n406), .O(n1078));
  nor2   g0763(.a(G55), .b(G18), .O(n1079));
  nor2   g0764(.a(n1079), .b(n1078), .O(n1080));
  inv1   g0765(.a(n1080), .O(n1081));
  nor2   g0766(.a(n1081), .b(n1077), .O(n1082));
  inv1   g0767(.a(n1077), .O(n1083));
  nor2   g0768(.a(n1080), .b(n1083), .O(n1084));
  nor2   g0769(.a(n1084), .b(n1082), .O(n1085));
  inv1   g0770(.a(n1085), .O(n1086));
  nor2   g0771(.a(n1086), .b(n1074), .O(n1087));
  inv1   g0772(.a(n1087), .O(n1088));
  nor2   g0773(.a(n1088), .b(n999), .O(n1089));
  nor2   g0774(.a(n1089), .b(n985), .O(n1090));
  inv1   g0775(.a(n1090), .O(n1091));
  inv1   g0776(.a(G187), .O(n1092));
  nor2   g0777(.a(n1092), .b(n406), .O(n1093));
  nor2   g0778(.a(n1093), .b(n624), .O(n1094));
  nor2   g0779(.a(n644), .b(n406), .O(n1095));
  nor2   g0780(.a(G77), .b(G18), .O(n1096));
  nor2   g0781(.a(n1096), .b(n1095), .O(n1097));
  inv1   g0782(.a(n1097), .O(n1098));
  nor2   g0783(.a(n1098), .b(n1094), .O(n1099));
  inv1   g0784(.a(n1082), .O(n1100));
  nor2   g0785(.a(n1100), .b(n995), .O(n1101));
  nor2   g0786(.a(n1101), .b(n1099), .O(n1102));
  inv1   g0787(.a(n1102), .O(n1103));
  nor2   g0788(.a(n1103), .b(n1091), .O(n1104));
  inv1   g0789(.a(G193), .O(n1105));
  nor2   g0790(.a(n1105), .b(n406), .O(n1106));
  nor2   g0791(.a(n1106), .b(n581), .O(n1107));
  inv1   g0792(.a(n1107), .O(n1108));
  nor2   g0793(.a(n584), .b(n406), .O(n1109));
  nor2   g0794(.a(G80), .b(G18), .O(n1110));
  nor2   g0795(.a(n1110), .b(n1109), .O(n1111));
  nor2   g0796(.a(n1111), .b(n1108), .O(n1112));
  inv1   g0797(.a(n1111), .O(n1113));
  nor2   g0798(.a(n1113), .b(n1107), .O(n1114));
  nor2   g0799(.a(n1114), .b(n1112), .O(n1115));
  inv1   g0800(.a(n1115), .O(n1116));
  inv1   g0801(.a(G194), .O(n1117));
  nor2   g0802(.a(n1117), .b(n406), .O(n1118));
  nor2   g0803(.a(n1118), .b(n592), .O(n1119));
  nor2   g0804(.a(n595), .b(n406), .O(n1120));
  nor2   g0805(.a(G81), .b(G18), .O(n1121));
  nor2   g0806(.a(n1121), .b(n1120), .O(n1122));
  inv1   g0807(.a(n1122), .O(n1123));
  nor2   g0808(.a(n1123), .b(n1119), .O(n1124));
  inv1   g0809(.a(n1119), .O(n1125));
  nor2   g0810(.a(n1122), .b(n1125), .O(n1126));
  nor2   g0811(.a(n1126), .b(n1124), .O(n1127));
  inv1   g0812(.a(n1127), .O(n1128));
  nor2   g0813(.a(n1128), .b(n1116), .O(n1129));
  inv1   g0814(.a(n1129), .O(n1130));
  inv1   g0815(.a(G196), .O(n1131));
  nor2   g0816(.a(n1131), .b(n406), .O(n1132));
  nor2   g0817(.a(n1132), .b(n611), .O(n1133));
  nor2   g0818(.a(n628), .b(n406), .O(n1134));
  nor2   g0819(.a(G78), .b(G18), .O(n1135));
  nor2   g0820(.a(n1135), .b(n1134), .O(n1136));
  inv1   g0821(.a(n1136), .O(n1137));
  nor2   g0822(.a(n1137), .b(n1133), .O(n1138));
  inv1   g0823(.a(G195), .O(n1139));
  nor2   g0824(.a(n1139), .b(n406), .O(n1140));
  nor2   g0825(.a(n1140), .b(n605), .O(n1141));
  inv1   g0826(.a(n1141), .O(n1142));
  nor2   g0827(.a(n615), .b(n406), .O(n1143));
  nor2   g0828(.a(G59), .b(G18), .O(n1144));
  nor2   g0829(.a(n1144), .b(n1143), .O(n1145));
  nor2   g0830(.a(n1145), .b(n1142), .O(n1146));
  nor2   g0831(.a(n1146), .b(n1138), .O(n1147));
  inv1   g0832(.a(n1147), .O(n1148));
  inv1   g0833(.a(n1133), .O(n1149));
  nor2   g0834(.a(n1136), .b(n1149), .O(n1150));
  inv1   g0835(.a(n1145), .O(n1151));
  nor2   g0836(.a(n1151), .b(n1141), .O(n1152));
  nor2   g0837(.a(n1152), .b(n1150), .O(n1153));
  inv1   g0838(.a(n1153), .O(n1154));
  nor2   g0839(.a(n1154), .b(n1148), .O(n1155));
  inv1   g0840(.a(n1155), .O(n1156));
  nor2   g0841(.a(n1156), .b(n1130), .O(n1157));
  inv1   g0842(.a(n1157), .O(n1158));
  inv1   g0843(.a(n1094), .O(n1159));
  nor2   g0844(.a(n1097), .b(n1159), .O(n1160));
  nor2   g0845(.a(n1160), .b(n1158), .O(n1161));
  inv1   g0846(.a(n1161), .O(n1162));
  nor2   g0847(.a(n1162), .b(n1104), .O(n1163));
  inv1   g0848(.a(n1138), .O(n1164));
  nor2   g0849(.a(n1146), .b(n1164), .O(n1165));
  nor2   g0850(.a(n1165), .b(n1152), .O(n1166));
  nor2   g0851(.a(n1166), .b(n1130), .O(n1167));
  inv1   g0852(.a(n1124), .O(n1168));
  nor2   g0853(.a(n1168), .b(n1112), .O(n1169));
  nor2   g0854(.a(n1169), .b(n1114), .O(n1170));
  inv1   g0855(.a(n1170), .O(n1171));
  nor2   g0856(.a(n1171), .b(n1167), .O(n1172));
  inv1   g0857(.a(n1172), .O(n1173));
  nor2   g0858(.a(n1173), .b(n1163), .O(n1174));
  nor2   g0859(.a(n1174), .b(n977), .O(n1175));
  inv1   g0860(.a(n947), .O(n1176));
  nor2   g0861(.a(n961), .b(n1176), .O(n1177));
  nor2   g0862(.a(n1177), .b(n963), .O(n1178));
  inv1   g0863(.a(n1178), .O(n1179));
  nor2   g0864(.a(n1179), .b(n1175), .O(n1180));
  inv1   g0865(.a(n1180), .O(n1181));
  nor2   g0866(.a(n1181), .b(n970), .O(n1182));
  nor2   g0867(.a(G174), .b(n406), .O(n1183));
  nor2   g0868(.a(n1183), .b(n405), .O(n1184));
  nor2   g0869(.a(n467), .b(n406), .O(n1185));
  nor2   g0870(.a(G109), .b(G18), .O(n1186));
  nor2   g0871(.a(n1186), .b(n1185), .O(n1187));
  nor2   g0872(.a(n1187), .b(n1184), .O(n1188));
  inv1   g0873(.a(n1184), .O(n1189));
  inv1   g0874(.a(n1187), .O(n1190));
  nor2   g0875(.a(n1190), .b(n1189), .O(n1191));
  nor2   g0876(.a(n1191), .b(n1188), .O(n1192));
  inv1   g0877(.a(n1192), .O(n1193));
  nor2   g0878(.a(G173), .b(n406), .O(n1194));
  nor2   g0879(.a(n1194), .b(n405), .O(n1195));
  nor2   g0880(.a(n471), .b(n406), .O(n1196));
  nor2   g0881(.a(G110), .b(G18), .O(n1197));
  nor2   g0882(.a(n1197), .b(n1196), .O(n1198));
  nor2   g0883(.a(n1198), .b(n1195), .O(n1199));
  inv1   g0884(.a(n1195), .O(n1200));
  inv1   g0885(.a(n1198), .O(n1201));
  nor2   g0886(.a(n1201), .b(n1200), .O(n1202));
  nor2   g0887(.a(n1202), .b(n1199), .O(n1203));
  inv1   g0888(.a(n1203), .O(n1204));
  nor2   g0889(.a(n1204), .b(n1193), .O(n1205));
  inv1   g0890(.a(n1205), .O(n1206));
  nor2   g0891(.a(G176), .b(n406), .O(n1207));
  nor2   g0892(.a(n1207), .b(n405), .O(n1208));
  nor2   g0893(.a(n493), .b(n406), .O(n1209));
  nor2   g0894(.a(G63), .b(G18), .O(n1210));
  nor2   g0895(.a(n1210), .b(n1209), .O(n1211));
  nor2   g0896(.a(n1211), .b(n1208), .O(n1212));
  nor2   g0897(.a(G175), .b(n406), .O(n1213));
  nor2   g0898(.a(n1213), .b(n405), .O(n1214));
  nor2   g0899(.a(n489), .b(n406), .O(n1215));
  nor2   g0900(.a(G86), .b(G18), .O(n1216));
  nor2   g0901(.a(n1216), .b(n1215), .O(n1217));
  nor2   g0902(.a(n1217), .b(n1214), .O(n1218));
  nor2   g0903(.a(n1218), .b(n1212), .O(n1219));
  inv1   g0904(.a(n1219), .O(n1220));
  inv1   g0905(.a(n1208), .O(n1221));
  inv1   g0906(.a(n1211), .O(n1222));
  nor2   g0907(.a(n1222), .b(n1221), .O(n1223));
  inv1   g0908(.a(n1214), .O(n1224));
  inv1   g0909(.a(n1217), .O(n1225));
  nor2   g0910(.a(n1225), .b(n1224), .O(n1226));
  nor2   g0911(.a(n1226), .b(n1223), .O(n1227));
  inv1   g0912(.a(n1227), .O(n1228));
  nor2   g0913(.a(n1228), .b(n1220), .O(n1229));
  inv1   g0914(.a(n1229), .O(n1230));
  nor2   g0915(.a(n1230), .b(n1206), .O(n1231));
  inv1   g0916(.a(n1231), .O(n1232));
  inv1   g0917(.a(G171), .O(n1233));
  nor2   g0918(.a(n1233), .b(n406), .O(n1234));
  nor2   g0919(.a(n1234), .b(n533), .O(n1235));
  nor2   g0920(.a(n825), .b(n406), .O(n1236));
  nor2   g0921(.a(G65), .b(G18), .O(n1237));
  nor2   g0922(.a(n1237), .b(n1236), .O(n1238));
  inv1   g0923(.a(n1238), .O(n1239));
  nor2   g0924(.a(n1239), .b(n1235), .O(n1240));
  inv1   g0925(.a(n1235), .O(n1241));
  nor2   g0926(.a(n1238), .b(n1241), .O(n1242));
  nor2   g0927(.a(n1242), .b(n1240), .O(n1243));
  inv1   g0928(.a(n1243), .O(n1244));
  nor2   g0929(.a(G177), .b(n406), .O(n1245));
  nor2   g0930(.a(n1245), .b(n405), .O(n1246));
  nor2   g0931(.a(n499), .b(n406), .O(n1247));
  nor2   g0932(.a(G64), .b(G18), .O(n1248));
  nor2   g0933(.a(n1248), .b(n1247), .O(n1249));
  nor2   g0934(.a(n1249), .b(n1246), .O(n1250));
  inv1   g0935(.a(n1246), .O(n1251));
  inv1   g0936(.a(n1249), .O(n1252));
  nor2   g0937(.a(n1252), .b(n1251), .O(n1253));
  nor2   g0938(.a(n1253), .b(n1250), .O(n1254));
  inv1   g0939(.a(n1254), .O(n1255));
  inv1   g0940(.a(G178), .O(n1256));
  nor2   g0941(.a(n1256), .b(n406), .O(n1257));
  nor2   g0942(.a(n1257), .b(n504), .O(n1258));
  nor2   g0943(.a(n509), .b(n406), .O(n1259));
  nor2   g0944(.a(G85), .b(G18), .O(n1260));
  nor2   g0945(.a(n1260), .b(n1259), .O(n1261));
  inv1   g0946(.a(n1261), .O(n1262));
  nor2   g0947(.a(n1262), .b(n1258), .O(n1263));
  inv1   g0948(.a(n1258), .O(n1264));
  nor2   g0949(.a(n1261), .b(n1264), .O(n1265));
  nor2   g0950(.a(n1265), .b(n1263), .O(n1266));
  inv1   g0951(.a(n1266), .O(n1267));
  nor2   g0952(.a(n1267), .b(n1255), .O(n1268));
  inv1   g0953(.a(n1268), .O(n1269));
  inv1   g0954(.a(G179), .O(n1270));
  nor2   g0955(.a(n1270), .b(n406), .O(n1271));
  nor2   g0956(.a(n1271), .b(n518), .O(n1272));
  inv1   g0957(.a(n1272), .O(n1273));
  nor2   g0958(.a(n516), .b(n406), .O(n1274));
  nor2   g0959(.a(G84), .b(G18), .O(n1275));
  nor2   g0960(.a(n1275), .b(n1274), .O(n1276));
  nor2   g0961(.a(n1276), .b(n1273), .O(n1277));
  inv1   g0962(.a(n1276), .O(n1278));
  nor2   g0963(.a(n1278), .b(n1272), .O(n1279));
  nor2   g0964(.a(n1279), .b(n1277), .O(n1280));
  inv1   g0965(.a(n1280), .O(n1281));
  inv1   g0966(.a(G180), .O(n1282));
  nor2   g0967(.a(n1282), .b(n406), .O(n1283));
  nor2   g0968(.a(n1283), .b(n526), .O(n1284));
  nor2   g0969(.a(n524), .b(n406), .O(n1285));
  nor2   g0970(.a(G83), .b(G18), .O(n1286));
  nor2   g0971(.a(n1286), .b(n1285), .O(n1287));
  inv1   g0972(.a(n1287), .O(n1288));
  nor2   g0973(.a(n1288), .b(n1284), .O(n1289));
  inv1   g0974(.a(n1284), .O(n1290));
  nor2   g0975(.a(n1287), .b(n1290), .O(n1291));
  nor2   g0976(.a(n1291), .b(n1289), .O(n1292));
  inv1   g0977(.a(n1292), .O(n1293));
  nor2   g0978(.a(n1293), .b(n1281), .O(n1294));
  inv1   g0979(.a(n1294), .O(n1295));
  nor2   g0980(.a(n1295), .b(n1269), .O(n1296));
  inv1   g0981(.a(n1296), .O(n1297));
  nor2   g0982(.a(n1297), .b(n1244), .O(n1298));
  inv1   g0983(.a(n1298), .O(n1299));
  nor2   g0984(.a(n1299), .b(n1232), .O(n1300));
  inv1   g0985(.a(n1300), .O(n1301));
  nor2   g0986(.a(n1301), .b(n1182), .O(n1302));
  inv1   g0987(.a(n1191), .O(n1303));
  nor2   g0988(.a(n1199), .b(n1303), .O(n1304));
  nor2   g0989(.a(n1304), .b(n1202), .O(n1305));
  inv1   g0990(.a(n1305), .O(n1306));
  inv1   g0991(.a(n1240), .O(n1307));
  nor2   g0992(.a(n1295), .b(n1307), .O(n1308));
  inv1   g0993(.a(n1289), .O(n1309));
  nor2   g0994(.a(n1309), .b(n1277), .O(n1310));
  nor2   g0995(.a(n1310), .b(n1279), .O(n1311));
  inv1   g0996(.a(n1311), .O(n1312));
  nor2   g0997(.a(n1312), .b(n1308), .O(n1313));
  nor2   g0998(.a(n1313), .b(n1269), .O(n1314));
  inv1   g0999(.a(n1263), .O(n1315));
  nor2   g1000(.a(n1315), .b(n1250), .O(n1316));
  nor2   g1001(.a(n1316), .b(n1253), .O(n1317));
  inv1   g1002(.a(n1317), .O(n1318));
  nor2   g1003(.a(n1318), .b(n1314), .O(n1319));
  nor2   g1004(.a(n1319), .b(n1232), .O(n1320));
  nor2   g1005(.a(n1227), .b(n1206), .O(n1321));
  inv1   g1006(.a(n1321), .O(n1322));
  nor2   g1007(.a(n1322), .b(n1218), .O(n1323));
  nor2   g1008(.a(n1323), .b(n1320), .O(n1324));
  inv1   g1009(.a(n1324), .O(n1325));
  nor2   g1010(.a(n1325), .b(n1306), .O(n1326));
  inv1   g1011(.a(n1326), .O(n1327));
  nor2   g1012(.a(n1327), .b(n1302), .O(n1328));
  inv1   g1013(.a(n405), .O(n1329));
  nor2   g1014(.a(n914), .b(n1329), .O(n1330));
  nor2   g1015(.a(n1330), .b(n916), .O(n1331));
  inv1   g1016(.a(n1331), .O(n1332));
  nor2   g1017(.a(n911), .b(n886), .O(n1333));
  inv1   g1018(.a(n1333), .O(n1334));
  inv1   g1019(.a(n874), .O(n1335));
  inv1   g1020(.a(n877), .O(n1336));
  nor2   g1021(.a(n1336), .b(n1335), .O(n1337));
  nor2   g1022(.a(n1337), .b(n878), .O(n1338));
  inv1   g1023(.a(n1338), .O(n1339));
  nor2   g1024(.a(n1339), .b(n1334), .O(n1340));
  inv1   g1025(.a(n1340), .O(n1341));
  nor2   g1026(.a(n1341), .b(n910), .O(n1342));
  inv1   g1027(.a(n1342), .O(n1343));
  nor2   g1028(.a(n1343), .b(n1332), .O(n1344));
  inv1   g1029(.a(n1344), .O(n1345));
  nor2   g1030(.a(n1345), .b(n1328), .O(n1346));
  nor2   g1031(.a(G2204), .b(G1455), .O(n1347));
  inv1   g1032(.a(n1347), .O(n1348));
  nor2   g1033(.a(n1348), .b(n387), .O(n1349));
  nor2   g1034(.a(n1349), .b(n385), .O(n1350));
  inv1   g1035(.a(n905), .O(n1351));
  nor2   g1036(.a(n1351), .b(n895), .O(n1352));
  nor2   g1037(.a(n1352), .b(n894), .O(n1353));
  nor2   g1038(.a(n1353), .b(n1341), .O(n1354));
  nor2   g1039(.a(n1354), .b(n1337), .O(n1355));
  inv1   g1040(.a(n1355), .O(n1356));
  nor2   g1041(.a(n1356), .b(n1350), .O(n1357));
  inv1   g1042(.a(n1357), .O(n1358));
  nor2   g1043(.a(n1358), .b(n1346), .O(n1359));
  inv1   g1044(.a(n1359), .O(n1360));
  nor2   g1045(.a(n1360), .b(n922), .O(n1361));
  nor2   g1046(.a(n1361), .b(n872), .O(G258));
  nor2   g1047(.a(n382), .b(n375), .O(n1363));
  nor2   g1048(.a(n1363), .b(n726), .O(n1364));
  nor2   g1049(.a(n1364), .b(n714), .O(n1365));
  nor2   g1050(.a(n1365), .b(n693), .O(n1366));
  nor2   g1051(.a(n1366), .b(n690), .O(n1367));
  inv1   g1052(.a(n1367), .O(n1368));
  nor2   g1053(.a(n1368), .b(n684), .O(n1369));
  nor2   g1054(.a(n1367), .b(n683), .O(n1370));
  nor2   g1055(.a(n1370), .b(n1369), .O(n1371));
  inv1   g1056(.a(n1371), .O(G388));
  nor2   g1057(.a(n1365), .b(n694), .O(n1373));
  inv1   g1058(.a(n1365), .O(n1374));
  nor2   g1059(.a(n1374), .b(n695), .O(n1375));
  nor2   g1060(.a(n1375), .b(n1373), .O(n1376));
  inv1   g1061(.a(n1376), .O(G391));
  nor2   g1062(.a(n712), .b(n375), .O(n1378));
  nor2   g1063(.a(n1378), .b(n722), .O(n1379));
  inv1   g1064(.a(n382), .O(n1380));
  nor2   g1065(.a(n724), .b(n1380), .O(n1381));
  nor2   g1066(.a(n1381), .b(n1379), .O(n1382));
  inv1   g1067(.a(n1382), .O(n1383));
  nor2   g1068(.a(n1383), .b(n719), .O(n1384));
  nor2   g1069(.a(n1382), .b(n718), .O(n1385));
  nor2   g1070(.a(n1385), .b(n1384), .O(n1386));
  inv1   g1071(.a(n1386), .O(G394));
  inv1   g1072(.a(n1363), .O(n1388));
  nor2   g1073(.a(n1388), .b(n723), .O(n1389));
  nor2   g1074(.a(n1363), .b(n724), .O(n1390));
  nor2   g1075(.a(n1390), .b(n1389), .O(G397));
  inv1   g1076(.a(n741), .O(n1392));
  inv1   g1077(.a(n778), .O(n1393));
  nor2   g1078(.a(n1393), .b(n1392), .O(n1394));
  nor2   g1079(.a(n673), .b(n665), .O(n1395));
  nor2   g1080(.a(n1395), .b(n660), .O(n1396));
  nor2   g1081(.a(n1396), .b(n766), .O(n1397));
  nor2   g1082(.a(n1397), .b(n763), .O(n1398));
  inv1   g1083(.a(n1398), .O(n1399));
  nor2   g1084(.a(n1399), .b(n741), .O(n1400));
  nor2   g1085(.a(n1400), .b(n1394), .O(n1401));
  inv1   g1086(.a(n1401), .O(n1402));
  nor2   g1087(.a(n1402), .b(n756), .O(n1403));
  nor2   g1088(.a(n1401), .b(n757), .O(n1404));
  nor2   g1089(.a(n1404), .b(n1403), .O(n1405));
  inv1   g1090(.a(n1405), .O(G376));
  inv1   g1091(.a(n776), .O(n1407));
  nor2   g1092(.a(n1407), .b(n1392), .O(n1408));
  nor2   g1093(.a(n1408), .b(n1396), .O(n1409));
  inv1   g1094(.a(n1409), .O(n1410));
  nor2   g1095(.a(n1410), .b(n767), .O(n1411));
  nor2   g1096(.a(n1409), .b(n768), .O(n1412));
  nor2   g1097(.a(n1412), .b(n1411), .O(n1413));
  inv1   g1098(.a(n1413), .O(G379));
  nor2   g1099(.a(n746), .b(n742), .O(n1415));
  inv1   g1100(.a(n1415), .O(n1416));
  nor2   g1101(.a(n1416), .b(n665), .O(n1417));
  nor2   g1102(.a(n1415), .b(n664), .O(n1418));
  nor2   g1103(.a(n1418), .b(n1417), .O(n1419));
  inv1   g1104(.a(n1419), .O(G382));
  nor2   g1105(.a(n746), .b(n673), .O(n1421));
  nor2   g1106(.a(n1421), .b(n1392), .O(n1422));
  inv1   g1107(.a(n1421), .O(n1423));
  nor2   g1108(.a(n1423), .b(n741), .O(n1424));
  nor2   g1109(.a(n1424), .b(n1422), .O(G385));
  inv1   g1110(.a(n485), .O(n1426));
  nor2   g1111(.a(n1426), .b(n483), .O(n1427));
  inv1   g1112(.a(n481), .O(n1428));
  nor2   g1113(.a(n487), .b(n1428), .O(n1429));
  nor2   g1114(.a(n1429), .b(n1427), .O(n1430));
  inv1   g1115(.a(n1430), .O(n1431));
  nor2   g1116(.a(n510), .b(n497), .O(n1432));
  nor2   g1117(.a(n507), .b(n496), .O(n1433));
  nor2   g1118(.a(n1433), .b(n1432), .O(n1434));
  nor2   g1119(.a(n1434), .b(n1431), .O(n1435));
  inv1   g1120(.a(n1434), .O(n1436));
  nor2   g1121(.a(n1436), .b(n1430), .O(n1437));
  nor2   g1122(.a(n1437), .b(n1435), .O(n1438));
  nor2   g1123(.a(n530), .b(n522), .O(n1439));
  nor2   g1124(.a(n529), .b(n521), .O(n1440));
  nor2   g1125(.a(n1440), .b(n1439), .O(n1441));
  inv1   g1126(.a(n1441), .O(n1442));
  inv1   g1127(.a(n472), .O(n1443));
  nor2   g1128(.a(n1443), .b(n465), .O(n1444));
  inv1   g1129(.a(n463), .O(n1445));
  nor2   g1130(.a(n475), .b(n1445), .O(n1446));
  nor2   g1131(.a(n1446), .b(n1444), .O(n1447));
  inv1   g1132(.a(n1447), .O(n1448));
  inv1   g1133(.a(G141), .O(n1449));
  nor2   g1134(.a(n1449), .b(G18), .O(n1450));
  inv1   g1135(.a(G161), .O(n1451));
  nor2   g1136(.a(n1451), .b(n406), .O(n1452));
  nor2   g1137(.a(n1452), .b(n1450), .O(n1453));
  nor2   g1138(.a(n1453), .b(n826), .O(n1454));
  inv1   g1139(.a(n1453), .O(n1455));
  nor2   g1140(.a(n1455), .b(n536), .O(n1456));
  nor2   g1141(.a(n1456), .b(n1454), .O(n1457));
  inv1   g1142(.a(n1457), .O(n1458));
  nor2   g1143(.a(n1458), .b(n1448), .O(n1459));
  nor2   g1144(.a(n1457), .b(n1447), .O(n1460));
  nor2   g1145(.a(n1460), .b(n1459), .O(n1461));
  nor2   g1146(.a(n1461), .b(n1442), .O(n1462));
  inv1   g1147(.a(n1461), .O(n1463));
  nor2   g1148(.a(n1463), .b(n1441), .O(n1464));
  nor2   g1149(.a(n1464), .b(n1462), .O(n1465));
  inv1   g1150(.a(n1465), .O(n1466));
  nor2   g1151(.a(n1466), .b(n1438), .O(n1467));
  inv1   g1152(.a(n1438), .O(n1468));
  nor2   g1153(.a(n1465), .b(n1468), .O(n1469));
  nor2   g1154(.a(n1469), .b(n1467), .O(n1470));
  nor2   g1155(.a(n765), .b(n754), .O(n1471));
  nor2   g1156(.a(n762), .b(n751), .O(n1472));
  nor2   g1157(.a(n1472), .b(n1471), .O(n1473));
  inv1   g1158(.a(n1473), .O(n1474));
  nor2   g1159(.a(n671), .b(n662), .O(n1475));
  nor2   g1160(.a(n672), .b(n659), .O(n1476));
  nor2   g1161(.a(n1476), .b(n1475), .O(n1477));
  nor2   g1162(.a(n721), .b(n704), .O(n1478));
  nor2   g1163(.a(n711), .b(n703), .O(n1479));
  nor2   g1164(.a(n1479), .b(n1478), .O(n1480));
  inv1   g1165(.a(n1480), .O(n1481));
  nor2   g1166(.a(n1481), .b(n1477), .O(n1482));
  inv1   g1167(.a(n1477), .O(n1483));
  nor2   g1168(.a(n1480), .b(n1483), .O(n1484));
  nor2   g1169(.a(n1484), .b(n1482), .O(n1485));
  nor2   g1170(.a(n1485), .b(n1474), .O(n1486));
  inv1   g1171(.a(n1485), .O(n1487));
  nor2   g1172(.a(n1487), .b(n1473), .O(n1488));
  nor2   g1173(.a(n1488), .b(n1486), .O(n1489));
  inv1   g1174(.a(G239), .O(n1490));
  nor2   g1175(.a(n1490), .b(n406), .O(n1491));
  inv1   g1176(.a(G44), .O(n1492));
  nor2   g1177(.a(n1492), .b(G18), .O(n1493));
  nor2   g1178(.a(n1493), .b(n1491), .O(n1494));
  inv1   g1179(.a(G229), .O(n1495));
  nor2   g1180(.a(n1495), .b(n406), .O(n1496));
  nor2   g1181(.a(n1496), .b(n373), .O(n1497));
  inv1   g1182(.a(n1497), .O(n1498));
  nor2   g1183(.a(n1498), .b(n1494), .O(n1499));
  inv1   g1184(.a(n1494), .O(n1500));
  nor2   g1185(.a(n1497), .b(n1500), .O(n1501));
  nor2   g1186(.a(n1501), .b(n1499), .O(n1502));
  inv1   g1187(.a(n1502), .O(n1503));
  nor2   g1188(.a(n692), .b(n681), .O(n1504));
  nor2   g1189(.a(n689), .b(n678), .O(n1505));
  nor2   g1190(.a(n1505), .b(n1504), .O(n1506));
  nor2   g1191(.a(n1506), .b(n1503), .O(n1507));
  inv1   g1192(.a(n1506), .O(n1508));
  nor2   g1193(.a(n1508), .b(n1502), .O(n1509));
  nor2   g1194(.a(n1509), .b(n1507), .O(n1510));
  nor2   g1195(.a(n1510), .b(n1489), .O(n1511));
  inv1   g1196(.a(n1489), .O(n1512));
  inv1   g1197(.a(n1510), .O(n1513));
  nor2   g1198(.a(n1513), .b(n1512), .O(n1514));
  nor2   g1199(.a(n1514), .b(n1511), .O(n1515));
  nor2   g1200(.a(n1515), .b(n1470), .O(n1516));
  inv1   g1201(.a(n1516), .O(n1517));
  nor2   g1202(.a(n596), .b(n585), .O(n1518));
  nor2   g1203(.a(n593), .b(n582), .O(n1519));
  nor2   g1204(.a(n1519), .b(n1518), .O(n1520));
  inv1   g1205(.a(G227), .O(n1521));
  nor2   g1206(.a(n1521), .b(n406), .O(n1522));
  inv1   g1207(.a(G115), .O(n1523));
  nor2   g1208(.a(n1523), .b(G18), .O(n1524));
  nor2   g1209(.a(n1524), .b(n1522), .O(n1525));
  inv1   g1210(.a(n1525), .O(n1526));
  nor2   g1211(.a(n1526), .b(n645), .O(n1527));
  nor2   g1212(.a(n1525), .b(n625), .O(n1528));
  nor2   g1213(.a(n1528), .b(n1527), .O(n1529));
  inv1   g1214(.a(n1529), .O(n1530));
  nor2   g1215(.a(n629), .b(n616), .O(n1531));
  nor2   g1216(.a(n612), .b(n606), .O(n1532));
  nor2   g1217(.a(n1532), .b(n1531), .O(n1533));
  nor2   g1218(.a(n1533), .b(n1530), .O(n1534));
  inv1   g1219(.a(n1533), .O(n1535));
  nor2   g1220(.a(n1535), .b(n1529), .O(n1536));
  nor2   g1221(.a(n1536), .b(n1534), .O(n1537));
  nor2   g1222(.a(n1537), .b(n1520), .O(n1538));
  inv1   g1223(.a(n1520), .O(n1539));
  inv1   g1224(.a(n1537), .O(n1540));
  nor2   g1225(.a(n1540), .b(n1539), .O(n1541));
  nor2   g1226(.a(n1541), .b(n1538), .O(n1542));
  nor2   g1227(.a(n806), .b(n796), .O(n1543));
  nor2   g1228(.a(n805), .b(n793), .O(n1544));
  nor2   g1229(.a(n1544), .b(n1543), .O(n1545));
  nor2   g1230(.a(n572), .b(n558), .O(n1546));
  nor2   g1231(.a(n569), .b(n561), .O(n1547));
  nor2   g1232(.a(n1547), .b(n1546), .O(n1548));
  inv1   g1233(.a(n1548), .O(n1549));
  nor2   g1234(.a(n1549), .b(n1545), .O(n1550));
  inv1   g1235(.a(n1545), .O(n1551));
  nor2   g1236(.a(n1548), .b(n1551), .O(n1552));
  nor2   g1237(.a(n1552), .b(n1550), .O(n1553));
  inv1   g1238(.a(n1553), .O(n1554));
  nor2   g1239(.a(n1554), .b(n1542), .O(n1555));
  inv1   g1240(.a(n1542), .O(n1556));
  nor2   g1241(.a(n1553), .b(n1556), .O(n1557));
  nor2   g1242(.a(n1557), .b(n1555), .O(n1558));
  inv1   g1243(.a(n1558), .O(n1559));
  nor2   g1244(.a(n405), .b(n406), .O(n1560));
  inv1   g1245(.a(n1560), .O(n1561));
  nor2   g1246(.a(G212), .b(G211), .O(n1562));
  inv1   g1247(.a(G211), .O(n1563));
  inv1   g1248(.a(G212), .O(n1564));
  nor2   g1249(.a(n1564), .b(n1563), .O(n1565));
  nor2   g1250(.a(n1565), .b(n1562), .O(n1566));
  inv1   g1251(.a(n1566), .O(n1567));
  nor2   g1252(.a(n1567), .b(G209), .O(n1568));
  inv1   g1253(.a(G209), .O(n1569));
  nor2   g1254(.a(n1566), .b(n1569), .O(n1570));
  nor2   g1255(.a(n1570), .b(n1568), .O(n1571));
  inv1   g1256(.a(n1571), .O(n1572));
  nor2   g1257(.a(n1572), .b(n1561), .O(n1573));
  inv1   g1258(.a(n444), .O(n1574));
  nor2   g1259(.a(n1574), .b(n436), .O(n1575));
  inv1   g1260(.a(n434), .O(n1576));
  nor2   g1261(.a(n446), .b(n1576), .O(n1577));
  nor2   g1262(.a(n1577), .b(n1575), .O(n1578));
  inv1   g1263(.a(n407), .O(n1579));
  nor2   g1264(.a(n415), .b(n1579), .O(n1580));
  inv1   g1265(.a(n413), .O(n1581));
  nor2   g1266(.a(n1581), .b(n409), .O(n1582));
  nor2   g1267(.a(n1582), .b(n1580), .O(n1583));
  inv1   g1268(.a(n1583), .O(n1584));
  nor2   g1269(.a(n1584), .b(n1578), .O(n1585));
  inv1   g1270(.a(n1578), .O(n1586));
  nor2   g1271(.a(n1583), .b(n1586), .O(n1587));
  nor2   g1272(.a(n1587), .b(n1585), .O(n1588));
  inv1   g1273(.a(n1588), .O(n1589));
  nor2   g1274(.a(n1589), .b(n1573), .O(n1590));
  inv1   g1275(.a(n1573), .O(n1591));
  nor2   g1276(.a(n1588), .b(n1591), .O(n1592));
  nor2   g1277(.a(n1592), .b(n1590), .O(n1593));
  nor2   g1278(.a(n1593), .b(n1559), .O(n1594));
  inv1   g1279(.a(n1594), .O(n1595));
  nor2   g1280(.a(n1595), .b(n1517), .O(n1596));
  inv1   g1281(.a(n1596), .O(G412));
  nor2   g1282(.a(n1217), .b(n1222), .O(n1598));
  nor2   g1283(.a(n1225), .b(n1211), .O(n1599));
  nor2   g1284(.a(n1599), .b(n1598), .O(n1600));
  inv1   g1285(.a(G2208), .O(n1601));
  nor2   g1286(.a(n1601), .b(n406), .O(n1602));
  nor2   g1287(.a(G82), .b(G18), .O(n1603));
  nor2   g1288(.a(n1603), .b(n1602), .O(n1604));
  inv1   g1289(.a(n1604), .O(n1605));
  nor2   g1290(.a(n1605), .b(n1239), .O(n1606));
  nor2   g1291(.a(n1604), .b(n1238), .O(n1607));
  nor2   g1292(.a(n1607), .b(n1606), .O(n1608));
  inv1   g1293(.a(n1608), .O(n1609));
  nor2   g1294(.a(n1609), .b(n1600), .O(n1610));
  inv1   g1295(.a(n1600), .O(n1611));
  nor2   g1296(.a(n1608), .b(n1611), .O(n1612));
  nor2   g1297(.a(n1612), .b(n1610), .O(n1613));
  nor2   g1298(.a(n1262), .b(n1252), .O(n1614));
  nor2   g1299(.a(n1261), .b(n1249), .O(n1615));
  nor2   g1300(.a(n1615), .b(n1614), .O(n1616));
  inv1   g1301(.a(n1616), .O(n1617));
  nor2   g1302(.a(n1288), .b(n1276), .O(n1618));
  nor2   g1303(.a(n1287), .b(n1278), .O(n1619));
  nor2   g1304(.a(n1619), .b(n1618), .O(n1620));
  inv1   g1305(.a(n1620), .O(n1621));
  nor2   g1306(.a(n1621), .b(n1617), .O(n1622));
  nor2   g1307(.a(n1620), .b(n1616), .O(n1623));
  nor2   g1308(.a(n1623), .b(n1622), .O(n1624));
  nor2   g1309(.a(n1201), .b(n1190), .O(n1625));
  nor2   g1310(.a(n1198), .b(n1187), .O(n1626));
  nor2   g1311(.a(n1626), .b(n1625), .O(n1627));
  inv1   g1312(.a(n1627), .O(n1628));
  nor2   g1313(.a(n1628), .b(n1624), .O(n1629));
  inv1   g1314(.a(n1624), .O(n1630));
  nor2   g1315(.a(n1627), .b(n1630), .O(n1631));
  nor2   g1316(.a(n1631), .b(n1629), .O(n1632));
  inv1   g1317(.a(n1632), .O(n1633));
  nor2   g1318(.a(n1633), .b(n1613), .O(n1634));
  inv1   g1319(.a(n1613), .O(n1635));
  nor2   g1320(.a(n1632), .b(n1635), .O(n1636));
  nor2   g1321(.a(n1636), .b(n1634), .O(n1637));
  nor2   g1322(.a(n904), .b(n893), .O(n1638));
  nor2   g1323(.a(n903), .b(n892), .O(n1639));
  nor2   g1324(.a(n1639), .b(n1638), .O(n1640));
  inv1   g1325(.a(n1640), .O(n1641));
  nor2   g1326(.a(n885), .b(n877), .O(n1642));
  nor2   g1327(.a(n884), .b(n1336), .O(n1643));
  nor2   g1328(.a(n1643), .b(n1642), .O(n1644));
  inv1   g1329(.a(n1644), .O(n1645));
  nor2   g1330(.a(n1645), .b(n1641), .O(n1646));
  nor2   g1331(.a(n1644), .b(n1640), .O(n1647));
  nor2   g1332(.a(n1647), .b(n1646), .O(n1648));
  inv1   g1333(.a(n1648), .O(n1649));
  nor2   g1334(.a(n393), .b(G1492), .O(n1650));
  nor2   g1335(.a(G1496), .b(n386), .O(n1651));
  nor2   g1336(.a(n1651), .b(n1650), .O(n1652));
  nor2   g1337(.a(n1652), .b(n406), .O(n1653));
  nor2   g1338(.a(n1347), .b(n871), .O(n1654));
  inv1   g1339(.a(n1654), .O(n1655));
  nor2   g1340(.a(n1655), .b(G18), .O(n1656));
  nor2   g1341(.a(n1656), .b(n1653), .O(n1657));
  inv1   g1342(.a(G1459), .O(n1658));
  nor2   g1343(.a(n1658), .b(n406), .O(n1659));
  nor2   g1344(.a(G114), .b(G18), .O(n1660));
  nor2   g1345(.a(n1660), .b(n1659), .O(n1661));
  inv1   g1346(.a(n1661), .O(n1662));
  nor2   g1347(.a(n1662), .b(n915), .O(n1663));
  nor2   g1348(.a(n1661), .b(n914), .O(n1664));
  nor2   g1349(.a(n1664), .b(n1663), .O(n1665));
  inv1   g1350(.a(n1665), .O(n1666));
  nor2   g1351(.a(n1666), .b(n1657), .O(n1667));
  inv1   g1352(.a(n1657), .O(n1668));
  nor2   g1353(.a(n1665), .b(n1668), .O(n1669));
  nor2   g1354(.a(n1669), .b(n1667), .O(n1670));
  inv1   g1355(.a(n1670), .O(n1671));
  nor2   g1356(.a(n1671), .b(n1649), .O(n1672));
  nor2   g1357(.a(n1670), .b(n1648), .O(n1673));
  nor2   g1358(.a(n1673), .b(n1672), .O(n1674));
  nor2   g1359(.a(n1674), .b(n1637), .O(n1675));
  inv1   g1360(.a(n1675), .O(n1676));
  nor2   g1361(.a(n1000), .b(n984), .O(n1677));
  nor2   g1362(.a(n992), .b(n983), .O(n1678));
  nor2   g1363(.a(n1678), .b(n1677), .O(n1679));
  nor2   g1364(.a(n376), .b(n406), .O(n1680));
  nor2   g1365(.a(n1680), .b(n1028), .O(n1681));
  inv1   g1366(.a(n1681), .O(n1682));
  inv1   g1367(.a(G3698), .O(n1683));
  nor2   g1368(.a(n1683), .b(n406), .O(n1684));
  nor2   g1369(.a(G69), .b(G18), .O(n1685));
  nor2   g1370(.a(n1685), .b(n1684), .O(n1686));
  inv1   g1371(.a(n1686), .O(n1687));
  nor2   g1372(.a(n1687), .b(n1682), .O(n1688));
  nor2   g1373(.a(n1686), .b(n1681), .O(n1689));
  nor2   g1374(.a(n1689), .b(n1688), .O(n1690));
  inv1   g1375(.a(n1690), .O(n1691));
  nor2   g1376(.a(n1691), .b(n1679), .O(n1692));
  inv1   g1377(.a(n1679), .O(n1693));
  nor2   g1378(.a(n1690), .b(n1693), .O(n1694));
  nor2   g1379(.a(n1694), .b(n1692), .O(n1695));
  nor2   g1380(.a(n1062), .b(n1060), .O(n1696));
  nor2   g1381(.a(n1053), .b(n1016), .O(n1697));
  nor2   g1382(.a(n1697), .b(n1696), .O(n1698));
  inv1   g1383(.a(n1698), .O(n1699));
  nor2   g1384(.a(n1039), .b(n1042), .O(n1700));
  nor2   g1385(.a(n1040), .b(n1025), .O(n1701));
  nor2   g1386(.a(n1701), .b(n1700), .O(n1702));
  inv1   g1387(.a(n1702), .O(n1703));
  nor2   g1388(.a(n1703), .b(n1699), .O(n1704));
  nor2   g1389(.a(n1702), .b(n1698), .O(n1705));
  nor2   g1390(.a(n1705), .b(n1704), .O(n1706));
  nor2   g1391(.a(n1080), .b(n1008), .O(n1707));
  nor2   g1392(.a(n1081), .b(n1007), .O(n1708));
  nor2   g1393(.a(n1708), .b(n1707), .O(n1709));
  inv1   g1394(.a(n1709), .O(n1710));
  nor2   g1395(.a(n1710), .b(n1706), .O(n1711));
  inv1   g1396(.a(n1706), .O(n1712));
  nor2   g1397(.a(n1709), .b(n1712), .O(n1713));
  nor2   g1398(.a(n1713), .b(n1711), .O(n1714));
  nor2   g1399(.a(n1714), .b(n1695), .O(n1715));
  inv1   g1400(.a(n1695), .O(n1716));
  inv1   g1401(.a(n1714), .O(n1717));
  nor2   g1402(.a(n1717), .b(n1716), .O(n1718));
  nor2   g1403(.a(n1718), .b(n1715), .O(n1719));
  inv1   g1404(.a(n1719), .O(n1720));
  nor2   g1405(.a(n1123), .b(n1113), .O(n1721));
  nor2   g1406(.a(n1122), .b(n1111), .O(n1722));
  nor2   g1407(.a(n1722), .b(n1721), .O(n1723));
  inv1   g1408(.a(G4393), .O(n1724));
  nor2   g1409(.a(n1724), .b(n406), .O(n1725));
  nor2   g1410(.a(G58), .b(G18), .O(n1726));
  nor2   g1411(.a(n1726), .b(n1725), .O(n1727));
  inv1   g1412(.a(n1727), .O(n1728));
  nor2   g1413(.a(n1728), .b(n1098), .O(n1729));
  nor2   g1414(.a(n1727), .b(n1097), .O(n1730));
  nor2   g1415(.a(n1730), .b(n1729), .O(n1731));
  inv1   g1416(.a(n1731), .O(n1732));
  nor2   g1417(.a(n1151), .b(n1137), .O(n1733));
  nor2   g1418(.a(n1145), .b(n1136), .O(n1734));
  nor2   g1419(.a(n1734), .b(n1733), .O(n1735));
  nor2   g1420(.a(n1735), .b(n1732), .O(n1736));
  inv1   g1421(.a(n1735), .O(n1737));
  nor2   g1422(.a(n1737), .b(n1731), .O(n1738));
  nor2   g1423(.a(n1738), .b(n1736), .O(n1739));
  nor2   g1424(.a(n1739), .b(n1723), .O(n1740));
  inv1   g1425(.a(n1723), .O(n1741));
  inv1   g1426(.a(n1739), .O(n1742));
  nor2   g1427(.a(n1742), .b(n1741), .O(n1743));
  nor2   g1428(.a(n1743), .b(n1740), .O(n1744));
  nor2   g1429(.a(n962), .b(n946), .O(n1745));
  nor2   g1430(.a(n960), .b(n945), .O(n1746));
  nor2   g1431(.a(n1746), .b(n1745), .O(n1747));
  nor2   g1432(.a(n937), .b(n928), .O(n1748));
  nor2   g1433(.a(n936), .b(n929), .O(n1749));
  nor2   g1434(.a(n1749), .b(n1748), .O(n1750));
  inv1   g1435(.a(n1750), .O(n1751));
  nor2   g1436(.a(n1751), .b(n1747), .O(n1752));
  inv1   g1437(.a(n1747), .O(n1753));
  nor2   g1438(.a(n1750), .b(n1753), .O(n1754));
  nor2   g1439(.a(n1754), .b(n1752), .O(n1755));
  inv1   g1440(.a(n1755), .O(n1756));
  nor2   g1441(.a(n1756), .b(n1744), .O(n1757));
  inv1   g1442(.a(n1744), .O(n1758));
  nor2   g1443(.a(n1755), .b(n1758), .O(n1759));
  nor2   g1444(.a(n1759), .b(n1757), .O(n1760));
  inv1   g1445(.a(n1760), .O(n1761));
  nor2   g1446(.a(n1761), .b(n1720), .O(n1762));
  inv1   g1447(.a(n1762), .O(n1763));
  nor2   g1448(.a(n1763), .b(n1676), .O(n1764));
  inv1   g1449(.a(n1764), .O(G414));
  nor2   g1450(.a(n957), .b(n948), .O(n1766));
  nor2   g1451(.a(n956), .b(n942), .O(n1767));
  nor2   g1452(.a(n1767), .b(n1766), .O(n1768));
  inv1   g1453(.a(n1768), .O(n1769));
  nor2   g1454(.a(n952), .b(n972), .O(n1770));
  nor2   g1455(.a(n933), .b(n925), .O(n1771));
  nor2   g1456(.a(n1771), .b(n1770), .O(n1772));
  nor2   g1457(.a(n1772), .b(n1769), .O(n1773));
  inv1   g1458(.a(n1772), .O(n1774));
  nor2   g1459(.a(n1774), .b(n1768), .O(n1775));
  nor2   g1460(.a(n1775), .b(n1773), .O(n1776));
  nor2   g1461(.a(n1125), .b(n1108), .O(n1777));
  nor2   g1462(.a(n1119), .b(n1107), .O(n1778));
  nor2   g1463(.a(n1778), .b(n1777), .O(n1779));
  inv1   g1464(.a(n1779), .O(n1780));
  inv1   g1465(.a(G197), .O(n1781));
  nor2   g1466(.a(n1781), .b(n406), .O(n1782));
  nor2   g1467(.a(n1782), .b(n1524), .O(n1783));
  inv1   g1468(.a(n1783), .O(n1784));
  nor2   g1469(.a(n1784), .b(n1094), .O(n1785));
  nor2   g1470(.a(n1783), .b(n1159), .O(n1786));
  nor2   g1471(.a(n1786), .b(n1785), .O(n1787));
  inv1   g1472(.a(n1787), .O(n1788));
  nor2   g1473(.a(n1788), .b(n1780), .O(n1789));
  nor2   g1474(.a(n1787), .b(n1779), .O(n1790));
  nor2   g1475(.a(n1790), .b(n1789), .O(n1791));
  nor2   g1476(.a(n1142), .b(n1149), .O(n1792));
  nor2   g1477(.a(n1141), .b(n1133), .O(n1793));
  nor2   g1478(.a(n1793), .b(n1792), .O(n1794));
  inv1   g1479(.a(n1794), .O(n1795));
  nor2   g1480(.a(n1795), .b(n1791), .O(n1796));
  inv1   g1481(.a(n1791), .O(n1797));
  nor2   g1482(.a(n1794), .b(n1797), .O(n1798));
  nor2   g1483(.a(n1798), .b(n1796), .O(n1799));
  inv1   g1484(.a(n1799), .O(n1800));
  nor2   g1485(.a(n1800), .b(n1776), .O(n1801));
  inv1   g1486(.a(n1776), .O(n1802));
  nor2   g1487(.a(n1799), .b(n1802), .O(n1803));
  nor2   g1488(.a(n1803), .b(n1801), .O(n1804));
  inv1   g1489(.a(n1804), .O(n1805));
  inv1   g1490(.a(n1213), .O(n1806));
  nor2   g1491(.a(n1806), .b(n1221), .O(n1807));
  inv1   g1492(.a(n1207), .O(n1808));
  nor2   g1493(.a(n1224), .b(n1808), .O(n1809));
  nor2   g1494(.a(n1809), .b(n1807), .O(n1810));
  inv1   g1495(.a(n1810), .O(n1811));
  inv1   g1496(.a(n1194), .O(n1812));
  nor2   g1497(.a(n1812), .b(n1189), .O(n1813));
  inv1   g1498(.a(n1183), .O(n1814));
  nor2   g1499(.a(n1200), .b(n1814), .O(n1815));
  nor2   g1500(.a(n1815), .b(n1813), .O(n1816));
  inv1   g1501(.a(n1816), .O(n1817));
  nor2   g1502(.a(n1817), .b(n1811), .O(n1818));
  nor2   g1503(.a(n1816), .b(n1810), .O(n1819));
  nor2   g1504(.a(n1819), .b(n1818), .O(n1820));
  inv1   g1505(.a(G181), .O(n1821));
  nor2   g1506(.a(n1821), .b(n406), .O(n1822));
  nor2   g1507(.a(n1822), .b(n1450), .O(n1823));
  inv1   g1508(.a(n1823), .O(n1824));
  nor2   g1509(.a(n1824), .b(n1235), .O(n1825));
  nor2   g1510(.a(n1823), .b(n1241), .O(n1826));
  nor2   g1511(.a(n1826), .b(n1825), .O(n1827));
  nor2   g1512(.a(n1258), .b(n1251), .O(n1828));
  nor2   g1513(.a(n1264), .b(n1246), .O(n1829));
  nor2   g1514(.a(n1829), .b(n1828), .O(n1830));
  inv1   g1515(.a(n1830), .O(n1831));
  nor2   g1516(.a(n1831), .b(n1827), .O(n1832));
  inv1   g1517(.a(n1827), .O(n1833));
  nor2   g1518(.a(n1830), .b(n1833), .O(n1834));
  nor2   g1519(.a(n1834), .b(n1832), .O(n1835));
  inv1   g1520(.a(n1835), .O(n1836));
  nor2   g1521(.a(n1290), .b(n1273), .O(n1837));
  nor2   g1522(.a(n1284), .b(n1272), .O(n1838));
  nor2   g1523(.a(n1838), .b(n1837), .O(n1839));
  nor2   g1524(.a(n1839), .b(n1836), .O(n1840));
  inv1   g1525(.a(n1839), .O(n1841));
  nor2   g1526(.a(n1841), .b(n1835), .O(n1842));
  nor2   g1527(.a(n1842), .b(n1840), .O(n1843));
  inv1   g1528(.a(n1843), .O(n1844));
  nor2   g1529(.a(n1844), .b(n1820), .O(n1845));
  inv1   g1530(.a(n1820), .O(n1846));
  nor2   g1531(.a(n1843), .b(n1846), .O(n1847));
  nor2   g1532(.a(n1847), .b(n1845), .O(n1848));
  inv1   g1533(.a(n1848), .O(n1849));
  nor2   g1534(.a(n1849), .b(n1805), .O(n1850));
  inv1   g1535(.a(n1850), .O(n1851));
  nor2   g1536(.a(G165), .b(G164), .O(n1852));
  inv1   g1537(.a(G164), .O(n1853));
  inv1   g1538(.a(G165), .O(n1854));
  nor2   g1539(.a(n1854), .b(n1853), .O(n1855));
  nor2   g1540(.a(n1855), .b(n1852), .O(n1856));
  inv1   g1541(.a(n1856), .O(n1857));
  nor2   g1542(.a(n1857), .b(G170), .O(n1858));
  inv1   g1543(.a(G170), .O(n1859));
  nor2   g1544(.a(n1856), .b(n1859), .O(n1860));
  nor2   g1545(.a(n1860), .b(n1858), .O(n1861));
  inv1   g1546(.a(n1861), .O(n1862));
  nor2   g1547(.a(n1862), .b(n1561), .O(n1863));
  inv1   g1548(.a(n1863), .O(n1864));
  inv1   g1549(.a(n887), .O(n1865));
  nor2   g1550(.a(n900), .b(n1865), .O(n1866));
  inv1   g1551(.a(n898), .O(n1867));
  nor2   g1552(.a(n1867), .b(n889), .O(n1868));
  nor2   g1553(.a(n1868), .b(n1866), .O(n1869));
  inv1   g1554(.a(n873), .O(n1870));
  nor2   g1555(.a(n881), .b(n1870), .O(n1871));
  inv1   g1556(.a(n879), .O(n1872));
  nor2   g1557(.a(n1872), .b(n1335), .O(n1873));
  nor2   g1558(.a(n1873), .b(n1871), .O(n1874));
  inv1   g1559(.a(n1874), .O(n1875));
  nor2   g1560(.a(n1875), .b(n1869), .O(n1876));
  inv1   g1561(.a(n1869), .O(n1877));
  nor2   g1562(.a(n1874), .b(n1877), .O(n1878));
  nor2   g1563(.a(n1878), .b(n1876), .O(n1879));
  inv1   g1564(.a(n1879), .O(n1880));
  nor2   g1565(.a(n1880), .b(n1864), .O(n1881));
  nor2   g1566(.a(n1879), .b(n1863), .O(n1882));
  nor2   g1567(.a(n1882), .b(n1881), .O(n1883));
  inv1   g1568(.a(n1883), .O(n1884));
  nor2   g1569(.a(n1077), .b(n1067), .O(n1885));
  nor2   g1570(.a(n1083), .b(n1004), .O(n1886));
  nor2   g1571(.a(n1886), .b(n1885), .O(n1887));
  inv1   g1572(.a(n1887), .O(n1888));
  inv1   g1573(.a(G198), .O(n1889));
  nor2   g1574(.a(n1889), .b(n406), .O(n1890));
  nor2   g1575(.a(n1890), .b(n373), .O(n1891));
  inv1   g1576(.a(n1891), .O(n1892));
  inv1   g1577(.a(G208), .O(n1893));
  nor2   g1578(.a(n1893), .b(n406), .O(n1894));
  nor2   g1579(.a(n1894), .b(n1493), .O(n1895));
  inv1   g1580(.a(n1895), .O(n1896));
  nor2   g1581(.a(n1896), .b(n1892), .O(n1897));
  nor2   g1582(.a(n1895), .b(n1891), .O(n1898));
  nor2   g1583(.a(n1898), .b(n1897), .O(n1899));
  nor2   g1584(.a(n1899), .b(n1888), .O(n1900));
  inv1   g1585(.a(n1899), .O(n1901));
  nor2   g1586(.a(n1901), .b(n1887), .O(n1902));
  nor2   g1587(.a(n1902), .b(n1900), .O(n1903));
  nor2   g1588(.a(n1050), .b(n1013), .O(n1904));
  nor2   g1589(.a(n1049), .b(n1012), .O(n1905));
  nor2   g1590(.a(n1905), .b(n1904), .O(n1906));
  inv1   g1591(.a(n1906), .O(n1907));
  nor2   g1592(.a(n1036), .b(n1022), .O(n1908));
  nor2   g1593(.a(n1055), .b(n1021), .O(n1909));
  nor2   g1594(.a(n1909), .b(n1908), .O(n1910));
  inv1   g1595(.a(n1910), .O(n1911));
  nor2   g1596(.a(n1911), .b(n1907), .O(n1912));
  nor2   g1597(.a(n1910), .b(n1906), .O(n1913));
  nor2   g1598(.a(n1913), .b(n1912), .O(n1914));
  nor2   g1599(.a(n989), .b(n994), .O(n1915));
  nor2   g1600(.a(n988), .b(n980), .O(n1916));
  nor2   g1601(.a(n1916), .b(n1915), .O(n1917));
  inv1   g1602(.a(n1917), .O(n1918));
  nor2   g1603(.a(n1918), .b(n1914), .O(n1919));
  inv1   g1604(.a(n1914), .O(n1920));
  nor2   g1605(.a(n1917), .b(n1920), .O(n1921));
  nor2   g1606(.a(n1921), .b(n1919), .O(n1922));
  inv1   g1607(.a(n1922), .O(n1923));
  nor2   g1608(.a(n1923), .b(n1903), .O(n1924));
  inv1   g1609(.a(n1903), .O(n1925));
  nor2   g1610(.a(n1922), .b(n1925), .O(n1926));
  nor2   g1611(.a(n1926), .b(n1924), .O(n1927));
  nor2   g1612(.a(n1927), .b(n1884), .O(n1928));
  inv1   g1613(.a(n1928), .O(n1929));
  nor2   g1614(.a(n1929), .b(n1851), .O(n1930));
  inv1   g1615(.a(n1930), .O(G416));
  nor2   g1616(.a(n829), .b(n820), .O(n1932));
  inv1   g1617(.a(n820), .O(n1933));
  nor2   g1618(.a(n828), .b(n1933), .O(n1934));
  nor2   g1619(.a(n1934), .b(n1932), .O(G295));
  inv1   g1620(.a(n853), .O(n1936));
  nor2   g1621(.a(n1936), .b(n461), .O(n1937));
  nor2   g1622(.a(n1937), .b(n854), .O(G324));
  inv1   g1623(.a(n1182), .O(G252));
  nor2   g1624(.a(n1932), .b(n537), .O(n1940));
  nor2   g1625(.a(n1940), .b(n824), .O(n1941));
  nor2   g1626(.a(n1941), .b(n543), .O(n1942));
  nor2   g1627(.a(n1942), .b(n523), .O(n1943));
  nor2   g1628(.a(n1943), .b(n508), .O(n1944));
  nor2   g1629(.a(n1944), .b(n511), .O(n1945));
  inv1   g1630(.a(n1945), .O(n1946));
  nor2   g1631(.a(n1946), .b(n501), .O(n1947));
  nor2   g1632(.a(n1945), .b(n502), .O(n1948));
  nor2   g1633(.a(n1948), .b(n1947), .O(n1949));
  inv1   g1634(.a(n1949), .O(G310));
  nor2   g1635(.a(n1943), .b(n512), .O(n1951));
  inv1   g1636(.a(n1943), .O(n1952));
  nor2   g1637(.a(n1952), .b(n513), .O(n1953));
  nor2   g1638(.a(n1953), .b(n1951), .O(G313));
  nor2   g1639(.a(n541), .b(n539), .O(n1955));
  inv1   g1640(.a(n1955), .O(n1956));
  nor2   g1641(.a(n831), .b(n820), .O(n1957));
  nor2   g1642(.a(n1957), .b(n1956), .O(n1958));
  inv1   g1643(.a(n1958), .O(n1959));
  nor2   g1644(.a(n1959), .b(n822), .O(n1960));
  nor2   g1645(.a(n1958), .b(n821), .O(n1961));
  nor2   g1646(.a(n1961), .b(n1960), .O(n1962));
  inv1   g1647(.a(n1962), .O(G316));
  inv1   g1648(.a(n1940), .O(n1964));
  nor2   g1649(.a(n1964), .b(n823), .O(n1965));
  nor2   g1650(.a(n1965), .b(n1941), .O(G319));
  nor2   g1651(.a(n456), .b(n416), .O(n1967));
  inv1   g1652(.a(n1967), .O(n1968));
  nor2   g1653(.a(n856), .b(n442), .O(n1969));
  nor2   g1654(.a(n1969), .b(n451), .O(n1970));
  nor2   g1655(.a(n1970), .b(n1968), .O(n1971));
  nor2   g1656(.a(n1971), .b(n424), .O(n1972));
  inv1   g1657(.a(n1972), .O(n1973));
  nor2   g1658(.a(n1973), .b(n421), .O(n1974));
  nor2   g1659(.a(n1972), .b(n422), .O(n1975));
  nor2   g1660(.a(n1975), .b(n1974), .O(n1976));
  inv1   g1661(.a(n1976), .O(G327));
  inv1   g1662(.a(n859), .O(n1978));
  nor2   g1663(.a(n1978), .b(n426), .O(n1979));
  nor2   g1664(.a(n859), .b(n425), .O(n1980));
  nor2   g1665(.a(n1980), .b(n1979), .O(n1981));
  inv1   g1666(.a(n1981), .O(G330));
  inv1   g1667(.a(n1969), .O(n1983));
  nor2   g1668(.a(n1983), .b(n437), .O(n1984));
  nor2   g1669(.a(n1984), .b(n450), .O(n1985));
  inv1   g1670(.a(n1984), .O(n1986));
  nor2   g1671(.a(n1986), .b(n451), .O(n1987));
  nor2   g1672(.a(n1987), .b(n1985), .O(n1988));
  inv1   g1673(.a(n1988), .O(G333));
  nor2   g1674(.a(n854), .b(n432), .O(n1990));
  inv1   g1675(.a(n1990), .O(n1991));
  nor2   g1676(.a(n1991), .b(n440), .O(n1992));
  nor2   g1677(.a(n1992), .b(n1983), .O(G336));
  nor2   g1678(.a(G416), .b(G408), .O(n1994));
  inv1   g1679(.a(n1994), .O(n1995));
  nor2   g1680(.a(n1995), .b(G410), .O(n1996));
  inv1   g1681(.a(n1996), .O(n1997));
  nor2   g1682(.a(G406), .b(G404), .O(n1998));
  inv1   g1683(.a(n1998), .O(n1999));
  nor2   g1684(.a(G414), .b(G412), .O(n2000));
  inv1   g1685(.a(n2000), .O(n2001));
  nor2   g1686(.a(n2001), .b(n1999), .O(n2002));
  inv1   g1687(.a(n2002), .O(n2003));
  nor2   g1688(.a(n2003), .b(n1997), .O(n2004));
  inv1   g1689(.a(n2004), .O(G418));
  nor2   g1690(.a(n494), .b(n492), .O(n2006));
  nor2   g1691(.a(n488), .b(n466), .O(n2007));
  inv1   g1692(.a(n2007), .O(n2008));
  nor2   g1693(.a(n2008), .b(n2006), .O(n2009));
  nor2   g1694(.a(n2009), .b(n468), .O(n2010));
  nor2   g1695(.a(n2010), .b(n837), .O(n2011));
  inv1   g1696(.a(n837), .O(n2012));
  nor2   g1697(.a(n850), .b(n2012), .O(n2013));
  nor2   g1698(.a(n2013), .b(n2011), .O(n2014));
  inv1   g1699(.a(n2014), .O(n2015));
  nor2   g1700(.a(n2015), .b(n478), .O(n2016));
  nor2   g1701(.a(n2014), .b(n477), .O(n2017));
  nor2   g1702(.a(n2017), .b(n2016), .O(G298));
  nor2   g1703(.a(n848), .b(n842), .O(n2019));
  nor2   g1704(.a(n2019), .b(n469), .O(n2020));
  inv1   g1705(.a(n2019), .O(n2021));
  nor2   g1706(.a(n2021), .b(n470), .O(n2022));
  nor2   g1707(.a(n2022), .b(n2020), .O(n2023));
  inv1   g1708(.a(n2023), .O(G301));
  nor2   g1709(.a(n491), .b(n484), .O(n2025));
  inv1   g1710(.a(n2025), .O(n2026));
  nor2   g1711(.a(n2026), .b(n838), .O(n2027));
  nor2   g1712(.a(n2027), .b(n840), .O(n2028));
  inv1   g1713(.a(n2028), .O(n2029));
  nor2   g1714(.a(n2029), .b(n846), .O(G304));
  nor2   g1715(.a(n494), .b(n484), .O(n2031));
  nor2   g1716(.a(n2031), .b(n2012), .O(n2032));
  inv1   g1717(.a(n2031), .O(n2033));
  nor2   g1718(.a(n2033), .b(n837), .O(n2034));
  nor2   g1719(.a(n2034), .b(n2032), .O(G307));
  nor2   g1720(.a(n782), .b(n648), .O(n2036));
  nor2   g1721(.a(n783), .b(n647), .O(n2037));
  nor2   g1722(.a(n2037), .b(n2036), .O(G344));
  nor2   g1723(.a(n389), .b(G38), .O(n2039));
  inv1   g1724(.a(n861), .O(n2040));
  nor2   g1725(.a(n863), .b(n2040), .O(n2041));
  nor2   g1726(.a(n2041), .b(n2039), .O(n2042));
  inv1   g1727(.a(n2042), .O(n2043));
  nor2   g1728(.a(n2043), .b(n399), .O(n2044));
  nor2   g1729(.a(n2042), .b(n400), .O(n2045));
  nor2   g1730(.a(n2045), .b(n2044), .O(n2046));
  inv1   g1731(.a(n2046), .O(G422));
  nor2   g1732(.a(n861), .b(n390), .O(n2048));
  inv1   g1733(.a(n2048), .O(n2049));
  nor2   g1734(.a(n2049), .b(n391), .O(n2050));
  inv1   g1735(.a(n2041), .O(n2051));
  nor2   g1736(.a(n2051), .b(n2039), .O(n2052));
  nor2   g1737(.a(n2052), .b(n2050), .O(n2053));
  inv1   g1738(.a(n2053), .O(G419));
  nor2   g1739(.a(n2036), .b(n626), .O(n2055));
  nor2   g1740(.a(n2055), .b(n650), .O(n2056));
  nor2   g1741(.a(n2056), .b(n620), .O(n2057));
  inv1   g1742(.a(n2057), .O(n2058));
  nor2   g1743(.a(n2058), .b(n594), .O(n2059));
  nor2   g1744(.a(n2059), .b(n597), .O(n2060));
  inv1   g1745(.a(n2060), .O(n2061));
  nor2   g1746(.a(n2061), .b(n587), .O(n2062));
  nor2   g1747(.a(n2060), .b(n588), .O(n2063));
  nor2   g1748(.a(n2063), .b(n2062), .O(n2064));
  inv1   g1749(.a(n2064), .O(G359));
  nor2   g1750(.a(n2058), .b(n598), .O(n2066));
  nor2   g1751(.a(n2057), .b(n599), .O(n2067));
  nor2   g1752(.a(n2067), .b(n2066), .O(G362));
  nor2   g1753(.a(n633), .b(n613), .O(n2069));
  inv1   g1754(.a(n2069), .O(n2070));
  nor2   g1755(.a(n648), .b(n632), .O(n2071));
  inv1   g1756(.a(n2071), .O(n2072));
  nor2   g1757(.a(n2072), .b(n782), .O(n2073));
  nor2   g1758(.a(n2073), .b(n2070), .O(n2074));
  inv1   g1759(.a(n2074), .O(n2075));
  nor2   g1760(.a(n2075), .b(n636), .O(n2076));
  nor2   g1761(.a(n2074), .b(n635), .O(n2077));
  nor2   g1762(.a(n2077), .b(n2076), .O(n2078));
  inv1   g1763(.a(n2078), .O(G365));
  inv1   g1764(.a(n2055), .O(n2080));
  nor2   g1765(.a(n2080), .b(n631), .O(n2081));
  nor2   g1766(.a(n2055), .b(n632), .O(n2082));
  nor2   g1767(.a(n2082), .b(n2081), .O(G368));
  inv1   g1768(.a(n817), .O(n2084));
  nor2   g1769(.a(n2084), .b(n785), .O(n2085));
  inv1   g1770(.a(n573), .O(n2086));
  nor2   g1771(.a(n2086), .b(n559), .O(n2087));
  nor2   g1772(.a(n797), .b(n562), .O(n2088));
  inv1   g1773(.a(n2088), .O(n2089));
  nor2   g1774(.a(n2089), .b(n2087), .O(n2090));
  nor2   g1775(.a(n2090), .b(n794), .O(n2091));
  nor2   g1776(.a(n2091), .b(n786), .O(n2092));
  nor2   g1777(.a(n2092), .b(n2085), .O(n2093));
  inv1   g1778(.a(n2093), .O(n2094));
  nor2   g1779(.a(n2094), .b(n810), .O(n2095));
  nor2   g1780(.a(n2093), .b(n809), .O(n2096));
  nor2   g1781(.a(n2096), .b(n2095), .O(n2097));
  inv1   g1782(.a(n2097), .O(G347));
  nor2   g1783(.a(n815), .b(n787), .O(n2099));
  inv1   g1784(.a(n2099), .O(n2100));
  nor2   g1785(.a(n2100), .b(n799), .O(n2101));
  nor2   g1786(.a(n2099), .b(n798), .O(n2102));
  nor2   g1787(.a(n2102), .b(n2101), .O(n2103));
  inv1   g1788(.a(n2103), .O(G350));
  nor2   g1789(.a(n785), .b(n570), .O(n2105));
  nor2   g1790(.a(n2105), .b(n573), .O(n2106));
  inv1   g1791(.a(n2106), .O(n2107));
  nor2   g1792(.a(n2107), .b(n564), .O(n2108));
  nor2   g1793(.a(n2106), .b(n563), .O(n2109));
  nor2   g1794(.a(n2109), .b(n2108), .O(G353));
  nor2   g1795(.a(n786), .b(n574), .O(n2111));
  nor2   g1796(.a(n785), .b(n575), .O(n2112));
  nor2   g1797(.a(n2112), .b(n2111), .O(n2113));
  inv1   g1798(.a(n2113), .O(G356));
  nor2   g1799(.a(n546), .b(n511), .O(n2115));
  nor2   g1800(.a(n545), .b(n508), .O(n2116));
  nor2   g1801(.a(n2116), .b(n2115), .O(n2117));
  inv1   g1802(.a(n2117), .O(n2118));
  nor2   g1803(.a(n828), .b(n823), .O(n2119));
  nor2   g1804(.a(n2119), .b(n830), .O(n2120));
  inv1   g1805(.a(n2120), .O(n2121));
  nor2   g1806(.a(n541), .b(n537), .O(n2122));
  nor2   g1807(.a(n2122), .b(n539), .O(n2123));
  inv1   g1808(.a(n2123), .O(n2124));
  nor2   g1809(.a(n2124), .b(n501), .O(n2125));
  nor2   g1810(.a(n2123), .b(n502), .O(n2126));
  nor2   g1811(.a(n2126), .b(n2125), .O(n2127));
  nor2   g1812(.a(n2127), .b(n2121), .O(n2128));
  inv1   g1813(.a(n2127), .O(n2129));
  nor2   g1814(.a(n2129), .b(n2120), .O(n2130));
  nor2   g1815(.a(n2130), .b(n2128), .O(n2131));
  inv1   g1816(.a(n2131), .O(n2132));
  nor2   g1817(.a(n2132), .b(n2118), .O(n2133));
  nor2   g1818(.a(n2131), .b(n2117), .O(n2134));
  nor2   g1819(.a(n2134), .b(n2133), .O(n2135));
  nor2   g1820(.a(n2135), .b(n1933), .O(n2136));
  nor2   g1821(.a(n833), .b(n513), .O(n2137));
  nor2   g1822(.a(n2115), .b(n508), .O(n2138));
  inv1   g1823(.a(n2138), .O(n2139));
  nor2   g1824(.a(n2139), .b(n2137), .O(n2140));
  inv1   g1825(.a(n2140), .O(n2141));
  nor2   g1826(.a(n2141), .b(n2120), .O(n2142));
  nor2   g1827(.a(n2140), .b(n2121), .O(n2143));
  nor2   g1828(.a(n2143), .b(n2142), .O(n2144));
  inv1   g1829(.a(n2144), .O(n2145));
  inv1   g1830(.a(n531), .O(n2146));
  nor2   g1831(.a(n827), .b(n2146), .O(n2147));
  inv1   g1832(.a(n541), .O(n2148));
  inv1   g1833(.a(n827), .O(n2149));
  nor2   g1834(.a(n2149), .b(n2148), .O(n2150));
  nor2   g1835(.a(n2150), .b(n2147), .O(n2151));
  inv1   g1836(.a(n2151), .O(n2152));
  nor2   g1837(.a(n832), .b(n545), .O(n2153));
  inv1   g1838(.a(n2153), .O(n2154));
  nor2   g1839(.a(n2154), .b(n502), .O(n2155));
  nor2   g1840(.a(n2153), .b(n501), .O(n2156));
  nor2   g1841(.a(n2156), .b(n2155), .O(n2157));
  nor2   g1842(.a(n2157), .b(n2152), .O(n2158));
  inv1   g1843(.a(n2157), .O(n2159));
  nor2   g1844(.a(n2159), .b(n2151), .O(n2160));
  nor2   g1845(.a(n2160), .b(n2158), .O(n2161));
  inv1   g1846(.a(n2161), .O(n2162));
  nor2   g1847(.a(n2162), .b(n2145), .O(n2163));
  nor2   g1848(.a(n2161), .b(n2144), .O(n2164));
  nor2   g1849(.a(n2164), .b(n2163), .O(n2165));
  nor2   g1850(.a(n2165), .b(n820), .O(n2166));
  nor2   g1851(.a(n2166), .b(n2136), .O(n2167));
  inv1   g1852(.a(n2167), .O(n2168));
  nor2   g1853(.a(n821), .b(n512), .O(n2169));
  nor2   g1854(.a(n822), .b(n513), .O(n2170));
  nor2   g1855(.a(n2170), .b(n2169), .O(n2171));
  nor2   g1856(.a(n834), .b(n553), .O(n2172));
  inv1   g1857(.a(n2172), .O(n2173));
  nor2   g1858(.a(n847), .b(n466), .O(n2174));
  nor2   g1859(.a(n2174), .b(n468), .O(n2175));
  inv1   g1860(.a(n2175), .O(n2176));
  nor2   g1861(.a(n847), .b(n494), .O(n2177));
  inv1   g1862(.a(n494), .O(n2178));
  nor2   g1863(.a(n2178), .b(n488), .O(n2179));
  nor2   g1864(.a(n2179), .b(n2177), .O(n2180));
  nor2   g1865(.a(n491), .b(n478), .O(n2181));
  nor2   g1866(.a(n492), .b(n477), .O(n2182));
  nor2   g1867(.a(n2182), .b(n2181), .O(n2183));
  inv1   g1868(.a(n2183), .O(n2184));
  nor2   g1869(.a(n2184), .b(n2180), .O(n2185));
  inv1   g1870(.a(n2180), .O(n2186));
  nor2   g1871(.a(n2183), .b(n2186), .O(n2187));
  nor2   g1872(.a(n2187), .b(n2185), .O(n2188));
  inv1   g1873(.a(n2188), .O(n2189));
  nor2   g1874(.a(n2189), .b(n2176), .O(n2190));
  nor2   g1875(.a(n2188), .b(n2175), .O(n2191));
  nor2   g1876(.a(n2191), .b(n2190), .O(n2192));
  inv1   g1877(.a(n2192), .O(n2193));
  nor2   g1878(.a(n2193), .b(n2173), .O(n2194));
  inv1   g1879(.a(n2010), .O(n2195));
  inv1   g1880(.a(n490), .O(n2196));
  nor2   g1881(.a(n2196), .b(n484), .O(n2197));
  nor2   g1882(.a(n2031), .b(n488), .O(n2198));
  nor2   g1883(.a(n2198), .b(n2025), .O(n2199));
  nor2   g1884(.a(n2199), .b(n2197), .O(n2200));
  nor2   g1885(.a(n477), .b(n469), .O(n2201));
  nor2   g1886(.a(n2201), .b(n479), .O(n2202));
  inv1   g1887(.a(n2202), .O(n2203));
  nor2   g1888(.a(n2203), .b(n2200), .O(n2204));
  inv1   g1889(.a(n2200), .O(n2205));
  nor2   g1890(.a(n2202), .b(n2205), .O(n2206));
  nor2   g1891(.a(n2206), .b(n2204), .O(n2207));
  inv1   g1892(.a(n2207), .O(n2208));
  nor2   g1893(.a(n2208), .b(n2195), .O(n2209));
  nor2   g1894(.a(n2207), .b(n2010), .O(n2210));
  nor2   g1895(.a(n2210), .b(n2209), .O(n2211));
  inv1   g1896(.a(n2211), .O(n2212));
  nor2   g1897(.a(n2212), .b(n2172), .O(n2213));
  nor2   g1898(.a(n2213), .b(n2194), .O(n2214));
  nor2   g1899(.a(n2214), .b(n820), .O(n2215));
  nor2   g1900(.a(n2212), .b(n552), .O(n2216));
  nor2   g1901(.a(n2193), .b(n553), .O(n2217));
  nor2   g1902(.a(n2217), .b(n2216), .O(n2218));
  nor2   g1903(.a(n2218), .b(n1933), .O(n2219));
  nor2   g1904(.a(n2219), .b(n2215), .O(n2220));
  inv1   g1905(.a(n2220), .O(n2221));
  nor2   g1906(.a(n2221), .b(n2171), .O(n2222));
  inv1   g1907(.a(n2171), .O(n2223));
  nor2   g1908(.a(n2220), .b(n2223), .O(n2224));
  nor2   g1909(.a(n2224), .b(n2222), .O(n2225));
  nor2   g1910(.a(n2225), .b(n2168), .O(n2226));
  inv1   g1911(.a(n2225), .O(n2227));
  nor2   g1912(.a(n2227), .b(n2167), .O(n2228));
  nor2   g1913(.a(n2228), .b(n2226), .O(G321));
  nor2   g1914(.a(n2048), .b(n391), .O(n2230));
  nor2   g1915(.a(n1968), .b(n452), .O(n2231));
  nor2   g1916(.a(n2231), .b(n424), .O(n2232));
  nor2   g1917(.a(n442), .b(n437), .O(n2233));
  nor2   g1918(.a(n2233), .b(n461), .O(n2234));
  nor2   g1919(.a(n462), .b(n437), .O(n2235));
  nor2   g1920(.a(n2235), .b(n2234), .O(n2236));
  nor2   g1921(.a(n2236), .b(n2232), .O(n2237));
  inv1   g1922(.a(n2232), .O(n2238));
  inv1   g1923(.a(n2236), .O(n2239));
  nor2   g1924(.a(n2239), .b(n2238), .O(n2240));
  nor2   g1925(.a(n2240), .b(n2237), .O(n2241));
  inv1   g1926(.a(n2241), .O(n2242));
  nor2   g1927(.a(n455), .b(n432), .O(n2243));
  nor2   g1928(.a(n458), .b(n433), .O(n2244));
  nor2   g1929(.a(n2244), .b(n2243), .O(n2245));
  inv1   g1930(.a(n2245), .O(n2246));
  nor2   g1931(.a(n441), .b(n421), .O(n2247));
  nor2   g1932(.a(n440), .b(n422), .O(n2248));
  nor2   g1933(.a(n2248), .b(n2247), .O(n2249));
  nor2   g1934(.a(n2249), .b(n2246), .O(n2250));
  inv1   g1935(.a(n2249), .O(n2251));
  nor2   g1936(.a(n2251), .b(n2245), .O(n2252));
  nor2   g1937(.a(n2252), .b(n2250), .O(n2253));
  inv1   g1938(.a(n2253), .O(n2254));
  nor2   g1939(.a(n2254), .b(n2242), .O(n2255));
  nor2   g1940(.a(n2253), .b(n2241), .O(n2256));
  nor2   g1941(.a(n2256), .b(n2255), .O(n2257));
  nor2   g1942(.a(n2257), .b(n1936), .O(n2258));
  nor2   g1943(.a(n460), .b(n441), .O(n2259));
  nor2   g1944(.a(n2259), .b(n437), .O(n2260));
  inv1   g1945(.a(n2260), .O(n2261));
  nor2   g1946(.a(n2261), .b(n421), .O(n2262));
  nor2   g1947(.a(n2260), .b(n422), .O(n2263));
  nor2   g1948(.a(n2263), .b(n2262), .O(n2264));
  inv1   g1949(.a(n2264), .O(n2265));
  inv1   g1950(.a(n2259), .O(n2266));
  nor2   g1951(.a(n2266), .b(n451), .O(n2267));
  nor2   g1952(.a(n460), .b(n456), .O(n2268));
  inv1   g1953(.a(n460), .O(n2269));
  nor2   g1954(.a(n2269), .b(n455), .O(n2270));
  nor2   g1955(.a(n2270), .b(n2268), .O(n2271));
  nor2   g1956(.a(n2271), .b(n2267), .O(n2272));
  inv1   g1957(.a(n2272), .O(n2273));
  nor2   g1958(.a(n2267), .b(n1968), .O(n2274));
  nor2   g1959(.a(n2274), .b(n424), .O(n2275));
  inv1   g1960(.a(n2275), .O(n2276));
  nor2   g1961(.a(n2266), .b(n432), .O(n2277));
  nor2   g1962(.a(n461), .b(n440), .O(n2278));
  nor2   g1963(.a(n2278), .b(n2277), .O(n2279));
  inv1   g1964(.a(n2279), .O(n2280));
  nor2   g1965(.a(n2280), .b(n2276), .O(n2281));
  nor2   g1966(.a(n2279), .b(n2275), .O(n2282));
  nor2   g1967(.a(n2282), .b(n2281), .O(n2283));
  nor2   g1968(.a(n2283), .b(n2273), .O(n2284));
  inv1   g1969(.a(n2283), .O(n2285));
  nor2   g1970(.a(n2285), .b(n2272), .O(n2286));
  nor2   g1971(.a(n2286), .b(n2284), .O(n2287));
  inv1   g1972(.a(n2287), .O(n2288));
  nor2   g1973(.a(n2288), .b(n2265), .O(n2289));
  nor2   g1974(.a(n2287), .b(n2264), .O(n2290));
  nor2   g1975(.a(n2290), .b(n2289), .O(n2291));
  nor2   g1976(.a(n2291), .b(n853), .O(n2292));
  nor2   g1977(.a(n2292), .b(n2258), .O(n2293));
  inv1   g1978(.a(n394), .O(n2294));
  nor2   g1979(.a(n426), .b(n2294), .O(n2295));
  nor2   g1980(.a(n425), .b(n394), .O(n2296));
  nor2   g1981(.a(n2296), .b(n2295), .O(n2297));
  nor2   g1982(.a(n2297), .b(n451), .O(n2298));
  inv1   g1983(.a(n2297), .O(n2299));
  nor2   g1984(.a(n2299), .b(n450), .O(n2300));
  nor2   g1985(.a(n2300), .b(n2298), .O(n2301));
  nor2   g1986(.a(n2301), .b(n2293), .O(n2302));
  inv1   g1987(.a(n2293), .O(n2303));
  inv1   g1988(.a(n2301), .O(n2304));
  nor2   g1989(.a(n2304), .b(n2303), .O(n2305));
  nor2   g1990(.a(n2305), .b(n2302), .O(n2306));
  nor2   g1991(.a(n2306), .b(n2230), .O(n2307));
  inv1   g1992(.a(n2230), .O(n2308));
  inv1   g1993(.a(n2306), .O(n2309));
  nor2   g1994(.a(n2309), .b(n2308), .O(n2310));
  nor2   g1995(.a(n2310), .b(n2307), .O(G338));
  inv1   g1996(.a(n815), .O(n2312));
  nor2   g1997(.a(n2312), .b(n794), .O(n2313));
  nor2   g1998(.a(n2313), .b(n797), .O(n2314));
  nor2   g1999(.a(n2312), .b(n573), .O(n2315));
  nor2   g2000(.a(n2315), .b(n2087), .O(n2316));
  inv1   g2001(.a(n2316), .O(n2317));
  nor2   g2002(.a(n810), .b(n564), .O(n2318));
  nor2   g2003(.a(n809), .b(n563), .O(n2319));
  nor2   g2004(.a(n2319), .b(n2318), .O(n2320));
  nor2   g2005(.a(n2320), .b(n2317), .O(n2321));
  inv1   g2006(.a(n2320), .O(n2322));
  nor2   g2007(.a(n2322), .b(n2316), .O(n2323));
  nor2   g2008(.a(n2323), .b(n2321), .O(n2324));
  nor2   g2009(.a(n2324), .b(n2314), .O(n2325));
  inv1   g2010(.a(n2314), .O(n2326));
  inv1   g2011(.a(n2324), .O(n2327));
  nor2   g2012(.a(n2327), .b(n2326), .O(n2328));
  nor2   g2013(.a(n2328), .b(n2325), .O(n2329));
  inv1   g2014(.a(n2329), .O(n2330));
  nor2   g2015(.a(n2330), .b(n643), .O(n2331));
  nor2   g2016(.a(n2316), .b(n563), .O(n2332));
  nor2   g2017(.a(n809), .b(n798), .O(n2333));
  nor2   g2018(.a(n2333), .b(n811), .O(n2334));
  inv1   g2019(.a(n2091), .O(n2335));
  nor2   g2020(.a(n2335), .b(n575), .O(n2336));
  nor2   g2021(.a(n2091), .b(n574), .O(n2337));
  nor2   g2022(.a(n2337), .b(n2336), .O(n2338));
  inv1   g2023(.a(n2338), .O(n2339));
  nor2   g2024(.a(n2339), .b(n2334), .O(n2340));
  inv1   g2025(.a(n2334), .O(n2341));
  nor2   g2026(.a(n2338), .b(n2341), .O(n2342));
  nor2   g2027(.a(n2342), .b(n2340), .O(n2343));
  nor2   g2028(.a(n2343), .b(n2332), .O(n2344));
  inv1   g2029(.a(n2332), .O(n2345));
  inv1   g2030(.a(n2343), .O(n2346));
  nor2   g2031(.a(n2346), .b(n2345), .O(n2347));
  nor2   g2032(.a(n2347), .b(n2344), .O(n2348));
  nor2   g2033(.a(n2348), .b(n642), .O(n2349));
  nor2   g2034(.a(n2349), .b(n2331), .O(n2350));
  inv1   g2035(.a(n2350), .O(n2351));
  nor2   g2036(.a(n2351), .b(n783), .O(n2352));
  nor2   g2037(.a(n2348), .b(n654), .O(n2353));
  inv1   g2038(.a(n654), .O(n2354));
  nor2   g2039(.a(n2330), .b(n2354), .O(n2355));
  nor2   g2040(.a(n2355), .b(n2353), .O(n2356));
  inv1   g2041(.a(n2356), .O(n2357));
  nor2   g2042(.a(n2357), .b(n782), .O(n2358));
  nor2   g2043(.a(n2358), .b(n2352), .O(n2359));
  inv1   g2044(.a(n646), .O(n2360));
  nor2   g2045(.a(n2360), .b(n614), .O(n2361));
  inv1   g2046(.a(n630), .O(n2362));
  nor2   g2047(.a(n646), .b(n2362), .O(n2363));
  nor2   g2048(.a(n2363), .b(n2361), .O(n2364));
  nor2   g2049(.a(n2360), .b(n631), .O(n2365));
  nor2   g2050(.a(n646), .b(n632), .O(n2366));
  nor2   g2051(.a(n2366), .b(n2365), .O(n2367));
  inv1   g2052(.a(n2367), .O(n2368));
  nor2   g2053(.a(n2368), .b(n626), .O(n2369));
  nor2   g2054(.a(n2369), .b(n633), .O(n2370));
  inv1   g2055(.a(n2370), .O(n2371));
  nor2   g2056(.a(n2371), .b(n587), .O(n2372));
  nor2   g2057(.a(n2370), .b(n588), .O(n2373));
  nor2   g2058(.a(n2373), .b(n2372), .O(n2374));
  inv1   g2059(.a(n2374), .O(n2375));
  nor2   g2060(.a(n2375), .b(n2364), .O(n2376));
  inv1   g2061(.a(n2364), .O(n2377));
  nor2   g2062(.a(n2374), .b(n2377), .O(n2378));
  nor2   g2063(.a(n2378), .b(n2376), .O(n2379));
  inv1   g2064(.a(n638), .O(n2380));
  nor2   g2065(.a(n651), .b(n2380), .O(n2381));
  inv1   g2066(.a(n2381), .O(n2382));
  nor2   g2067(.a(n652), .b(n599), .O(n2383));
  nor2   g2068(.a(n2380), .b(n594), .O(n2384));
  nor2   g2069(.a(n2384), .b(n597), .O(n2385));
  nor2   g2070(.a(n2385), .b(n2383), .O(n2386));
  inv1   g2071(.a(n2386), .O(n2387));
  nor2   g2072(.a(n2387), .b(n2382), .O(n2388));
  nor2   g2073(.a(n2386), .b(n2381), .O(n2389));
  nor2   g2074(.a(n2389), .b(n2388), .O(n2390));
  inv1   g2075(.a(n2390), .O(n2391));
  nor2   g2076(.a(n2391), .b(n2379), .O(n2392));
  inv1   g2077(.a(n2379), .O(n2393));
  nor2   g2078(.a(n2390), .b(n2393), .O(n2394));
  nor2   g2079(.a(n2394), .b(n2392), .O(n2395));
  nor2   g2080(.a(n2395), .b(n782), .O(n2396));
  inv1   g2081(.a(n2385), .O(n2397));
  nor2   g2082(.a(n2368), .b(n588), .O(n2398));
  nor2   g2083(.a(n2367), .b(n587), .O(n2399));
  nor2   g2084(.a(n2399), .b(n2398), .O(n2400));
  inv1   g2085(.a(n607), .O(n2401));
  nor2   g2086(.a(n2070), .b(n2401), .O(n2402));
  inv1   g2087(.a(n617), .O(n2403));
  nor2   g2088(.a(n2069), .b(n2403), .O(n2404));
  nor2   g2089(.a(n2404), .b(n2402), .O(n2405));
  inv1   g2090(.a(n2405), .O(n2406));
  nor2   g2091(.a(n2406), .b(n2400), .O(n2407));
  inv1   g2092(.a(n2400), .O(n2408));
  nor2   g2093(.a(n2405), .b(n2408), .O(n2409));
  nor2   g2094(.a(n2409), .b(n2407), .O(n2410));
  inv1   g2095(.a(n2410), .O(n2411));
  nor2   g2096(.a(n2411), .b(n2397), .O(n2412));
  nor2   g2097(.a(n2410), .b(n2385), .O(n2413));
  nor2   g2098(.a(n2413), .b(n2412), .O(n2414));
  nor2   g2099(.a(n2414), .b(n783), .O(n2415));
  nor2   g2100(.a(n2415), .b(n2396), .O(n2416));
  inv1   g2101(.a(n2416), .O(n2417));
  nor2   g2102(.a(n636), .b(n599), .O(n2418));
  nor2   g2103(.a(n635), .b(n598), .O(n2419));
  nor2   g2104(.a(n2419), .b(n2418), .O(n2420));
  nor2   g2105(.a(n2420), .b(n2417), .O(n2421));
  inv1   g2106(.a(n2420), .O(n2422));
  nor2   g2107(.a(n2422), .b(n2416), .O(n2423));
  nor2   g2108(.a(n2423), .b(n2421), .O(n2424));
  nor2   g2109(.a(n2424), .b(n2359), .O(n2425));
  inv1   g2110(.a(n2359), .O(n2426));
  inv1   g2111(.a(n2424), .O(n2427));
  nor2   g2112(.a(n2427), .b(n2426), .O(n2428));
  nor2   g2113(.a(n2428), .b(n2425), .O(n2429));
  inv1   g2114(.a(n2429), .O(G370));
  inv1   g2115(.a(n1396), .O(n2431));
  nor2   g2116(.a(n2431), .b(n766), .O(n2432));
  nor2   g2117(.a(n2432), .b(n763), .O(n2433));
  inv1   g2118(.a(n2433), .O(n2434));
  inv1   g2119(.a(n660), .O(n2435));
  nor2   g2120(.a(n746), .b(n2435), .O(n2436));
  inv1   g2121(.a(n673), .O(n2437));
  nor2   g2122(.a(n2437), .b(n663), .O(n2438));
  nor2   g2123(.a(n2438), .b(n746), .O(n2439));
  nor2   g2124(.a(n2439), .b(n660), .O(n2440));
  nor2   g2125(.a(n2440), .b(n2436), .O(n2441));
  inv1   g2126(.a(n2441), .O(n2442));
  nor2   g2127(.a(n2442), .b(n756), .O(n2443));
  nor2   g2128(.a(n2441), .b(n757), .O(n2444));
  nor2   g2129(.a(n2444), .b(n2443), .O(n2445));
  inv1   g2130(.a(n2445), .O(n2446));
  nor2   g2131(.a(n2446), .b(n2434), .O(n2447));
  nor2   g2132(.a(n2445), .b(n2433), .O(n2448));
  nor2   g2133(.a(n2448), .b(n2447), .O(n2449));
  nor2   g2134(.a(n2449), .b(n734), .O(n2450));
  nor2   g2135(.a(n776), .b(n763), .O(n2451));
  nor2   g2136(.a(n2451), .b(n766), .O(n2452));
  inv1   g2137(.a(n2452), .O(n2453));
  nor2   g2138(.a(n756), .b(n665), .O(n2454));
  nor2   g2139(.a(n757), .b(n664), .O(n2455));
  nor2   g2140(.a(n2455), .b(n2454), .O(n2456));
  inv1   g2141(.a(n2456), .O(n2457));
  nor2   g2142(.a(n1423), .b(n660), .O(n2458));
  inv1   g2143(.a(n663), .O(n2459));
  nor2   g2144(.a(n774), .b(n2459), .O(n2460));
  nor2   g2145(.a(n2460), .b(n2436), .O(n2461));
  nor2   g2146(.a(n2461), .b(n1421), .O(n2462));
  nor2   g2147(.a(n2462), .b(n2458), .O(n2463));
  inv1   g2148(.a(n2463), .O(n2464));
  nor2   g2149(.a(n2464), .b(n2457), .O(n2465));
  nor2   g2150(.a(n2463), .b(n2456), .O(n2466));
  nor2   g2151(.a(n2466), .b(n2465), .O(n2467));
  inv1   g2152(.a(n2467), .O(n2468));
  nor2   g2153(.a(n2468), .b(n2453), .O(n2469));
  nor2   g2154(.a(n2467), .b(n2452), .O(n2470));
  nor2   g2155(.a(n2470), .b(n2469), .O(n2471));
  nor2   g2156(.a(n2471), .b(n735), .O(n2472));
  nor2   g2157(.a(n2472), .b(G4526), .O(n2473));
  inv1   g2158(.a(n2473), .O(n2474));
  nor2   g2159(.a(n2474), .b(n2450), .O(n2475));
  nor2   g2160(.a(n738), .b(n735), .O(n2476));
  nor2   g2161(.a(n2476), .b(n2449), .O(n2477));
  inv1   g2162(.a(n2476), .O(n2478));
  nor2   g2163(.a(n2478), .b(n2471), .O(n2479));
  nor2   g2164(.a(n2479), .b(n371), .O(n2480));
  inv1   g2165(.a(n2480), .O(n2481));
  nor2   g2166(.a(n2481), .b(n2477), .O(n2482));
  nor2   g2167(.a(n2482), .b(n2475), .O(n2483));
  inv1   g2168(.a(n2483), .O(n2484));
  nor2   g2169(.a(n694), .b(n683), .O(n2485));
  nor2   g2170(.a(n2485), .b(n696), .O(n2486));
  nor2   g2171(.a(n2486), .b(n719), .O(n2487));
  inv1   g2172(.a(n2486), .O(n2488));
  nor2   g2173(.a(n2488), .b(n718), .O(n2489));
  nor2   g2174(.a(n2489), .b(n2487), .O(n2490));
  inv1   g2175(.a(n2490), .O(n2491));
  nor2   g2176(.a(n724), .b(n381), .O(n2492));
  nor2   g2177(.a(n723), .b(n380), .O(n2493));
  nor2   g2178(.a(n2493), .b(n2492), .O(n2494));
  inv1   g2179(.a(n2494), .O(n2495));
  nor2   g2180(.a(n727), .b(n714), .O(n2496));
  nor2   g2181(.a(n2496), .b(n693), .O(n2497));
  nor2   g2182(.a(n2497), .b(n690), .O(n2498));
  inv1   g2183(.a(n2498), .O(n2499));
  nor2   g2184(.a(n2499), .b(n2495), .O(n2500));
  nor2   g2185(.a(n2498), .b(n2494), .O(n2501));
  nor2   g2186(.a(n2501), .b(n2500), .O(n2502));
  inv1   g2187(.a(n2502), .O(n2503));
  nor2   g2188(.a(n714), .b(n375), .O(n2504));
  nor2   g2189(.a(n2496), .b(n717), .O(n2505));
  nor2   g2190(.a(n2505), .b(n2504), .O(n2506));
  inv1   g2191(.a(n2506), .O(n2507));
  nor2   g2192(.a(n2507), .b(n1379), .O(n2508));
  inv1   g2193(.a(n1379), .O(n2509));
  nor2   g2194(.a(n2506), .b(n2509), .O(n2510));
  nor2   g2195(.a(n2510), .b(n2508), .O(n2511));
  inv1   g2196(.a(n2511), .O(n2512));
  nor2   g2197(.a(n2512), .b(n2503), .O(n2513));
  nor2   g2198(.a(n2511), .b(n2502), .O(n2514));
  nor2   g2199(.a(n2514), .b(G4526), .O(n2515));
  inv1   g2200(.a(n2515), .O(n2516));
  nor2   g2201(.a(n2516), .b(n2513), .O(n2517));
  nor2   g2202(.a(n722), .b(n379), .O(n2518));
  inv1   g2203(.a(n379), .O(n2519));
  nor2   g2204(.a(n1379), .b(n2519), .O(n2520));
  nor2   g2205(.a(n2520), .b(n2518), .O(n2521));
  inv1   g2206(.a(n2521), .O(n2522));
  nor2   g2207(.a(n2522), .b(n2495), .O(n2523));
  nor2   g2208(.a(n2521), .b(n2494), .O(n2524));
  nor2   g2209(.a(n2524), .b(n2523), .O(n2525));
  inv1   g2210(.a(n2496), .O(n2526));
  nor2   g2211(.a(n2526), .b(n736), .O(n2527));
  nor2   g2212(.a(n2527), .b(n693), .O(n2528));
  inv1   g2213(.a(n2527), .O(n2529));
  nor2   g2214(.a(n2529), .b(n690), .O(n2530));
  nor2   g2215(.a(n2530), .b(n2528), .O(n2531));
  inv1   g2216(.a(n2531), .O(n2532));
  nor2   g2217(.a(n2532), .b(n2525), .O(n2533));
  inv1   g2218(.a(n2525), .O(n2534));
  nor2   g2219(.a(n2531), .b(n2534), .O(n2535));
  nor2   g2220(.a(n2535), .b(n2533), .O(n2536));
  inv1   g2221(.a(n2536), .O(n2537));
  nor2   g2222(.a(n2537), .b(n371), .O(n2538));
  nor2   g2223(.a(n2538), .b(n2517), .O(n2539));
  inv1   g2224(.a(n2539), .O(n2540));
  nor2   g2225(.a(n2540), .b(n2491), .O(n2541));
  nor2   g2226(.a(n2539), .b(n2490), .O(n2542));
  nor2   g2227(.a(n2542), .b(n2541), .O(n2543));
  inv1   g2228(.a(n2543), .O(n2544));
  nor2   g2229(.a(n2544), .b(n2484), .O(n2545));
  nor2   g2230(.a(n2543), .b(n2483), .O(n2546));
  nor2   g2231(.a(n2546), .b(n2545), .O(G399));
  buffer g2232(.a(ING339 ), .O(G339));
  buffer g2233(.a(G1), .O(G2));
  buffer g2234(.a(G1), .O(G3));
  buffer g2235(.a(G1459), .O(G450));
  buffer g2236(.a(G1469), .O(G448));
  buffer g2237(.a(G1480), .O(G444));
  buffer g2238(.a(G1486), .O(G442));
  buffer g2239(.a(G1492), .O(G440));
  buffer g2240(.a(G1496), .O(G438));
  buffer g2241(.a(G2208), .O(G496));
  buffer g2242(.a(G2218), .O(G494));
  buffer g2243(.a(G2224), .O(G492));
  buffer g2244(.a(G2230), .O(G490));
  buffer g2245(.a(G2236), .O(G488));
  buffer g2246(.a(G2239), .O(G486));
  buffer g2247(.a(G2247), .O(G484));
  buffer g2248(.a(G2253), .O(G482));
  buffer g2249(.a(G2256), .O(G480));
  buffer g2250(.a(G3698), .O(G560));
  buffer g2251(.a(G3701), .O(G542));
  buffer g2252(.a(G3705), .O(G558));
  buffer g2253(.a(G3711), .O(G556));
  buffer g2254(.a(G3717), .O(G554));
  buffer g2255(.a(G3723), .O(G552));
  buffer g2256(.a(G3729), .O(G550));
  buffer g2257(.a(G3737), .O(G548));
  buffer g2258(.a(G3743), .O(G546));
  buffer g2259(.a(G3749), .O(G544));
  buffer g2260(.a(G4393), .O(G540));
  buffer g2261(.a(G4400), .O(G538));
  buffer g2262(.a(G4405), .O(G536));
  buffer g2263(.a(G4410), .O(G534));
  buffer g2264(.a(G4415), .O(G532));
  buffer g2265(.a(G4420), .O(G530));
  buffer g2266(.a(G4427), .O(G528));
  buffer g2267(.a(G4432), .O(G526));
  buffer g2268(.a(G4437), .O(G524));
  buffer g2269(.a(G1462), .O(G436));
  buffer g2270(.a(G2211), .O(G478));
  buffer g2271(.a(G4394), .O(G522));
  buffer g2272(.a(G1), .O(G432));
  buffer g2273(.a(G106), .O(G446));
  inv1   g2274(.a(G15), .O(G286));
  inv1   g2275(.a(n360), .O(G289));
  inv1   g2276(.a(G15), .O(G341));
  inv1   g2277(.a(n366), .O(G281));
  buffer g2278(.a(G1), .O(G453));
  nor2   g2279(.a(n1361), .b(n872), .O(G264));
  inv1   g2280(.a(n867), .O(G270));
  nor2   g2281(.a(n1361), .b(n872), .O(G249));
  inv1   g2282(.a(n867), .O(G276));
  inv1   g2283(.a(n867), .O(G273));
  inv1   g2284(.a(n2046), .O(G469));
  inv1   g2285(.a(n2053), .O(G471));
endmodule


