// Benchmark "c6288_blif" written by ABC on Sun Mar 24 18:39:15 2019

module c6288_blif  ( 
    G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat,
    G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat,
    G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat,
    G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat,
    G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat  );
  input  G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat,
    G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat,
    G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat,
    G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat;
  output G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat;
  wire n65, n66, n68, n69, n70, n71, n72, n73, n74, n75, n76, n78, n79, n80,
    n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
    n95, n96, n97, n98, n100, n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n131, n132,
    n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
    n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
    n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467, n468, n469, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n575, n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n691,
    n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
    n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
    n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
    n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
    n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
    n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
    n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
    n812, n813, n814, n815, n816, n817, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
    n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
    n957, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
    n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
    n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
    n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
    n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
    n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
    n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
    n1105, n1106, n1107, n1108, n1109, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
    n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
    n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
    n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
    n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
    n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
    n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
    n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
    n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
    n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
    n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
    n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
    n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
    n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
    n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
    n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
    n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
    n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
    n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
    n1789, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
    n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
    n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
    n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
    n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
    n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
    n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
    n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
    n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
    n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
    n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
    n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
    n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
    n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
    n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
    n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
    n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
    n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
    n2222, n2223, n2224, n2225, n2226, n2228, n2229, n2230, n2231, n2232,
    n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
    n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
    n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
    n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
    n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
    n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
    n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348, n2350, n2351, n2352, n2353,
    n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
    n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
    n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
    n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
    n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
    n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
    n2454, n2455, n2456, n2457, n2458, n2460, n2461, n2462, n2463, n2464,
    n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
    n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
    n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
    n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
    n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
    n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
    n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
    n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
    n2555, n2556, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
    n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
    n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
    n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
    n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
    n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2644, n2645, n2646,
    n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
    n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
    n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
    n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
    n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
    n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
    n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
    n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
    n2778, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
    n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
    n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
    n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
    n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
    n2891, n2892, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
    n2902, n2903, n2905, n2906, n2907;
  inv1   g0000(.a(G1gat), .O(n65));
  inv1   g0001(.a(G273gat), .O(n66));
  nor2   g0002(.a(n66), .b(n65), .O(G545gat));
  inv1   g0003(.a(G18gat), .O(n68));
  nor2   g0004(.a(n66), .b(n68), .O(n69));
  inv1   g0005(.a(n69), .O(n70));
  inv1   g0006(.a(G290gat), .O(n71));
  nor2   g0007(.a(n71), .b(n65), .O(n72));
  nor2   g0008(.a(n72), .b(n70), .O(n73));
  inv1   g0009(.a(n72), .O(n74));
  nor2   g0010(.a(n74), .b(n69), .O(n75));
  nor2   g0011(.a(n75), .b(n73), .O(n76));
  inv1   g0012(.a(n76), .O(G1581gat));
  inv1   g0013(.a(G307gat), .O(n78));
  nor2   g0014(.a(n78), .b(n65), .O(n79));
  inv1   g0015(.a(G545gat), .O(n80));
  nor2   g0016(.a(n80), .b(G35gat), .O(n81));
  inv1   g0017(.a(G35gat), .O(n82));
  nor2   g0018(.a(n66), .b(n82), .O(n83));
  nor2   g0019(.a(n71), .b(n68), .O(n84));
  nor2   g0020(.a(n84), .b(n83), .O(n85));
  inv1   g0021(.a(n84), .O(n86));
  inv1   g0022(.a(n83), .O(n87));
  nor2   g0023(.a(n87), .b(G1gat), .O(n88));
  inv1   g0024(.a(n88), .O(n89));
  nor2   g0025(.a(n89), .b(n86), .O(n90));
  nor2   g0026(.a(n90), .b(n85), .O(n91));
  inv1   g0027(.a(n91), .O(n92));
  nor2   g0028(.a(n92), .b(n81), .O(n93));
  inv1   g0029(.a(n93), .O(n94));
  nor2   g0030(.a(n94), .b(n79), .O(n95));
  inv1   g0031(.a(n79), .O(n96));
  nor2   g0032(.a(n93), .b(n96), .O(n97));
  nor2   g0033(.a(n97), .b(n95), .O(n98));
  inv1   g0034(.a(n98), .O(G1901gat));
  inv1   g0035(.a(G324gat), .O(n100));
  nor2   g0036(.a(n100), .b(n65), .O(n101));
  nor2   g0037(.a(n95), .b(n92), .O(n102));
  nor2   g0038(.a(n78), .b(n68), .O(n103));
  inv1   g0039(.a(G52gat), .O(n104));
  nor2   g0040(.a(n66), .b(n104), .O(n105));
  inv1   g0041(.a(n105), .O(n106));
  nor2   g0042(.a(n71), .b(n82), .O(n107));
  inv1   g0043(.a(n107), .O(n108));
  nor2   g0044(.a(n108), .b(G18gat), .O(n109));
  nor2   g0045(.a(n109), .b(n106), .O(n110));
  nor2   g0046(.a(n108), .b(n105), .O(n111));
  inv1   g0047(.a(n111), .O(n112));
  nor2   g0048(.a(n112), .b(n69), .O(n113));
  nor2   g0049(.a(n113), .b(n110), .O(n114));
  nor2   g0050(.a(n114), .b(n103), .O(n115));
  inv1   g0051(.a(n103), .O(n116));
  inv1   g0052(.a(n114), .O(n117));
  nor2   g0053(.a(n117), .b(n116), .O(n118));
  nor2   g0054(.a(n118), .b(n115), .O(n119));
  inv1   g0055(.a(n119), .O(n120));
  nor2   g0056(.a(n120), .b(n102), .O(n121));
  inv1   g0057(.a(n102), .O(n122));
  nor2   g0058(.a(n119), .b(n122), .O(n123));
  nor2   g0059(.a(n123), .b(n121), .O(n124));
  inv1   g0060(.a(n124), .O(n125));
  nor2   g0061(.a(n125), .b(n101), .O(n126));
  inv1   g0062(.a(n101), .O(n127));
  nor2   g0063(.a(n124), .b(n127), .O(n128));
  nor2   g0064(.a(n128), .b(n126), .O(n129));
  inv1   g0065(.a(n129), .O(G2223gat));
  inv1   g0066(.a(G341gat), .O(n131));
  nor2   g0067(.a(n131), .b(n65), .O(n132));
  nor2   g0068(.a(n126), .b(n121), .O(n133));
  nor2   g0069(.a(n100), .b(n68), .O(n134));
  nor2   g0070(.a(n111), .b(n110), .O(n135));
  nor2   g0071(.a(n135), .b(n115), .O(n136));
  nor2   g0072(.a(n78), .b(n82), .O(n137));
  inv1   g0073(.a(G69gat), .O(n138));
  nor2   g0074(.a(n66), .b(n138), .O(n139));
  inv1   g0075(.a(n139), .O(n140));
  nor2   g0076(.a(n71), .b(n104), .O(n141));
  inv1   g0077(.a(n141), .O(n142));
  nor2   g0078(.a(n142), .b(G35gat), .O(n143));
  nor2   g0079(.a(n143), .b(n140), .O(n144));
  nor2   g0080(.a(n142), .b(n139), .O(n145));
  inv1   g0081(.a(n145), .O(n146));
  nor2   g0082(.a(n146), .b(n83), .O(n147));
  nor2   g0083(.a(n147), .b(n144), .O(n148));
  nor2   g0084(.a(n148), .b(n137), .O(n149));
  inv1   g0085(.a(n137), .O(n150));
  inv1   g0086(.a(n148), .O(n151));
  nor2   g0087(.a(n151), .b(n150), .O(n152));
  nor2   g0088(.a(n152), .b(n149), .O(n153));
  inv1   g0089(.a(n153), .O(n154));
  nor2   g0090(.a(n154), .b(n136), .O(n155));
  inv1   g0091(.a(n136), .O(n156));
  nor2   g0092(.a(n153), .b(n156), .O(n157));
  nor2   g0093(.a(n157), .b(n155), .O(n158));
  inv1   g0094(.a(n158), .O(n159));
  nor2   g0095(.a(n159), .b(n134), .O(n160));
  inv1   g0096(.a(n134), .O(n161));
  nor2   g0097(.a(n158), .b(n161), .O(n162));
  nor2   g0098(.a(n162), .b(n160), .O(n163));
  inv1   g0099(.a(n163), .O(n164));
  nor2   g0100(.a(n164), .b(n133), .O(n165));
  inv1   g0101(.a(n133), .O(n166));
  nor2   g0102(.a(n163), .b(n166), .O(n167));
  nor2   g0103(.a(n167), .b(n165), .O(n168));
  inv1   g0104(.a(n168), .O(n169));
  nor2   g0105(.a(n169), .b(n132), .O(n170));
  inv1   g0106(.a(n132), .O(n171));
  nor2   g0107(.a(n168), .b(n171), .O(n172));
  nor2   g0108(.a(n172), .b(n170), .O(n173));
  inv1   g0109(.a(n173), .O(G2548gat));
  inv1   g0110(.a(G358gat), .O(n175));
  nor2   g0111(.a(n175), .b(n65), .O(n176));
  nor2   g0112(.a(n170), .b(n165), .O(n177));
  nor2   g0113(.a(n131), .b(n68), .O(n178));
  nor2   g0114(.a(n160), .b(n155), .O(n179));
  nor2   g0115(.a(n100), .b(n82), .O(n180));
  nor2   g0116(.a(n145), .b(n144), .O(n181));
  nor2   g0117(.a(n181), .b(n149), .O(n182));
  nor2   g0118(.a(n78), .b(n104), .O(n183));
  inv1   g0119(.a(G86gat), .O(n184));
  nor2   g0120(.a(n66), .b(n184), .O(n185));
  inv1   g0121(.a(n185), .O(n186));
  nor2   g0122(.a(n71), .b(n138), .O(n187));
  inv1   g0123(.a(n187), .O(n188));
  nor2   g0124(.a(n188), .b(G52gat), .O(n189));
  nor2   g0125(.a(n189), .b(n186), .O(n190));
  nor2   g0126(.a(n188), .b(n185), .O(n191));
  inv1   g0127(.a(n191), .O(n192));
  nor2   g0128(.a(n192), .b(n105), .O(n193));
  nor2   g0129(.a(n193), .b(n190), .O(n194));
  nor2   g0130(.a(n194), .b(n183), .O(n195));
  inv1   g0131(.a(n183), .O(n196));
  inv1   g0132(.a(n194), .O(n197));
  nor2   g0133(.a(n197), .b(n196), .O(n198));
  nor2   g0134(.a(n198), .b(n195), .O(n199));
  inv1   g0135(.a(n199), .O(n200));
  nor2   g0136(.a(n200), .b(n182), .O(n201));
  inv1   g0137(.a(n182), .O(n202));
  nor2   g0138(.a(n199), .b(n202), .O(n203));
  nor2   g0139(.a(n203), .b(n201), .O(n204));
  inv1   g0140(.a(n204), .O(n205));
  nor2   g0141(.a(n205), .b(n180), .O(n206));
  inv1   g0142(.a(n180), .O(n207));
  nor2   g0143(.a(n204), .b(n207), .O(n208));
  nor2   g0144(.a(n208), .b(n206), .O(n209));
  inv1   g0145(.a(n209), .O(n210));
  nor2   g0146(.a(n210), .b(n179), .O(n211));
  inv1   g0147(.a(n179), .O(n212));
  nor2   g0148(.a(n209), .b(n212), .O(n213));
  nor2   g0149(.a(n213), .b(n211), .O(n214));
  inv1   g0150(.a(n214), .O(n215));
  nor2   g0151(.a(n215), .b(n178), .O(n216));
  inv1   g0152(.a(n178), .O(n217));
  nor2   g0153(.a(n214), .b(n217), .O(n218));
  nor2   g0154(.a(n218), .b(n216), .O(n219));
  inv1   g0155(.a(n219), .O(n220));
  nor2   g0156(.a(n220), .b(n177), .O(n221));
  inv1   g0157(.a(n177), .O(n222));
  nor2   g0158(.a(n219), .b(n222), .O(n223));
  nor2   g0159(.a(n223), .b(n221), .O(n224));
  inv1   g0160(.a(n224), .O(n225));
  nor2   g0161(.a(n225), .b(n176), .O(n226));
  inv1   g0162(.a(n176), .O(n227));
  nor2   g0163(.a(n224), .b(n227), .O(n228));
  nor2   g0164(.a(n228), .b(n226), .O(n229));
  inv1   g0165(.a(n229), .O(G2877gat));
  inv1   g0166(.a(G375gat), .O(n231));
  nor2   g0167(.a(n231), .b(n65), .O(n232));
  nor2   g0168(.a(n226), .b(n221), .O(n233));
  nor2   g0169(.a(n175), .b(n68), .O(n234));
  nor2   g0170(.a(n216), .b(n211), .O(n235));
  nor2   g0171(.a(n131), .b(n82), .O(n236));
  nor2   g0172(.a(n206), .b(n201), .O(n237));
  nor2   g0173(.a(n100), .b(n104), .O(n238));
  nor2   g0174(.a(n191), .b(n190), .O(n239));
  nor2   g0175(.a(n239), .b(n195), .O(n240));
  nor2   g0176(.a(n78), .b(n138), .O(n241));
  inv1   g0177(.a(G103gat), .O(n242));
  nor2   g0178(.a(n66), .b(n242), .O(n243));
  inv1   g0179(.a(n243), .O(n244));
  nor2   g0180(.a(n71), .b(n184), .O(n245));
  inv1   g0181(.a(n245), .O(n246));
  nor2   g0182(.a(n246), .b(G69gat), .O(n247));
  nor2   g0183(.a(n247), .b(n244), .O(n248));
  nor2   g0184(.a(n246), .b(n243), .O(n249));
  inv1   g0185(.a(n249), .O(n250));
  nor2   g0186(.a(n250), .b(n139), .O(n251));
  nor2   g0187(.a(n251), .b(n248), .O(n252));
  nor2   g0188(.a(n252), .b(n241), .O(n253));
  inv1   g0189(.a(n241), .O(n254));
  inv1   g0190(.a(n252), .O(n255));
  nor2   g0191(.a(n255), .b(n254), .O(n256));
  nor2   g0192(.a(n256), .b(n253), .O(n257));
  inv1   g0193(.a(n257), .O(n258));
  nor2   g0194(.a(n258), .b(n240), .O(n259));
  inv1   g0195(.a(n240), .O(n260));
  nor2   g0196(.a(n257), .b(n260), .O(n261));
  nor2   g0197(.a(n261), .b(n259), .O(n262));
  inv1   g0198(.a(n262), .O(n263));
  nor2   g0199(.a(n263), .b(n238), .O(n264));
  inv1   g0200(.a(n238), .O(n265));
  nor2   g0201(.a(n262), .b(n265), .O(n266));
  nor2   g0202(.a(n266), .b(n264), .O(n267));
  inv1   g0203(.a(n267), .O(n268));
  nor2   g0204(.a(n268), .b(n237), .O(n269));
  inv1   g0205(.a(n237), .O(n270));
  nor2   g0206(.a(n267), .b(n270), .O(n271));
  nor2   g0207(.a(n271), .b(n269), .O(n272));
  inv1   g0208(.a(n272), .O(n273));
  nor2   g0209(.a(n273), .b(n236), .O(n274));
  inv1   g0210(.a(n236), .O(n275));
  nor2   g0211(.a(n272), .b(n275), .O(n276));
  nor2   g0212(.a(n276), .b(n274), .O(n277));
  inv1   g0213(.a(n277), .O(n278));
  nor2   g0214(.a(n278), .b(n235), .O(n279));
  inv1   g0215(.a(n235), .O(n280));
  nor2   g0216(.a(n277), .b(n280), .O(n281));
  nor2   g0217(.a(n281), .b(n279), .O(n282));
  inv1   g0218(.a(n282), .O(n283));
  nor2   g0219(.a(n283), .b(n234), .O(n284));
  inv1   g0220(.a(n234), .O(n285));
  nor2   g0221(.a(n282), .b(n285), .O(n286));
  nor2   g0222(.a(n286), .b(n284), .O(n287));
  inv1   g0223(.a(n287), .O(n288));
  nor2   g0224(.a(n288), .b(n233), .O(n289));
  inv1   g0225(.a(n233), .O(n290));
  nor2   g0226(.a(n287), .b(n290), .O(n291));
  nor2   g0227(.a(n291), .b(n289), .O(n292));
  inv1   g0228(.a(n292), .O(n293));
  nor2   g0229(.a(n293), .b(n232), .O(n294));
  inv1   g0230(.a(n232), .O(n295));
  nor2   g0231(.a(n292), .b(n295), .O(n296));
  nor2   g0232(.a(n296), .b(n294), .O(n297));
  inv1   g0233(.a(n297), .O(G3211gat));
  inv1   g0234(.a(G392gat), .O(n299));
  nor2   g0235(.a(n299), .b(n65), .O(n300));
  nor2   g0236(.a(n294), .b(n289), .O(n301));
  nor2   g0237(.a(n231), .b(n68), .O(n302));
  nor2   g0238(.a(n284), .b(n279), .O(n303));
  nor2   g0239(.a(n175), .b(n82), .O(n304));
  nor2   g0240(.a(n274), .b(n269), .O(n305));
  nor2   g0241(.a(n131), .b(n104), .O(n306));
  nor2   g0242(.a(n264), .b(n259), .O(n307));
  nor2   g0243(.a(n100), .b(n138), .O(n308));
  nor2   g0244(.a(n249), .b(n248), .O(n309));
  nor2   g0245(.a(n309), .b(n253), .O(n310));
  nor2   g0246(.a(n78), .b(n184), .O(n311));
  inv1   g0247(.a(G120gat), .O(n312));
  nor2   g0248(.a(n66), .b(n312), .O(n313));
  inv1   g0249(.a(n313), .O(n314));
  nor2   g0250(.a(n71), .b(n242), .O(n315));
  inv1   g0251(.a(n315), .O(n316));
  nor2   g0252(.a(n316), .b(G86gat), .O(n317));
  nor2   g0253(.a(n317), .b(n314), .O(n318));
  nor2   g0254(.a(n316), .b(n313), .O(n319));
  inv1   g0255(.a(n319), .O(n320));
  nor2   g0256(.a(n320), .b(n185), .O(n321));
  nor2   g0257(.a(n321), .b(n318), .O(n322));
  nor2   g0258(.a(n322), .b(n311), .O(n323));
  inv1   g0259(.a(n311), .O(n324));
  inv1   g0260(.a(n322), .O(n325));
  nor2   g0261(.a(n325), .b(n324), .O(n326));
  nor2   g0262(.a(n326), .b(n323), .O(n327));
  inv1   g0263(.a(n327), .O(n328));
  nor2   g0264(.a(n328), .b(n310), .O(n329));
  inv1   g0265(.a(n310), .O(n330));
  nor2   g0266(.a(n327), .b(n330), .O(n331));
  nor2   g0267(.a(n331), .b(n329), .O(n332));
  inv1   g0268(.a(n332), .O(n333));
  nor2   g0269(.a(n333), .b(n308), .O(n334));
  inv1   g0270(.a(n308), .O(n335));
  nor2   g0271(.a(n332), .b(n335), .O(n336));
  nor2   g0272(.a(n336), .b(n334), .O(n337));
  inv1   g0273(.a(n337), .O(n338));
  nor2   g0274(.a(n338), .b(n307), .O(n339));
  inv1   g0275(.a(n307), .O(n340));
  nor2   g0276(.a(n337), .b(n340), .O(n341));
  nor2   g0277(.a(n341), .b(n339), .O(n342));
  inv1   g0278(.a(n342), .O(n343));
  nor2   g0279(.a(n343), .b(n306), .O(n344));
  inv1   g0280(.a(n306), .O(n345));
  nor2   g0281(.a(n342), .b(n345), .O(n346));
  nor2   g0282(.a(n346), .b(n344), .O(n347));
  inv1   g0283(.a(n347), .O(n348));
  nor2   g0284(.a(n348), .b(n305), .O(n349));
  inv1   g0285(.a(n305), .O(n350));
  nor2   g0286(.a(n347), .b(n350), .O(n351));
  nor2   g0287(.a(n351), .b(n349), .O(n352));
  inv1   g0288(.a(n352), .O(n353));
  nor2   g0289(.a(n353), .b(n304), .O(n354));
  inv1   g0290(.a(n304), .O(n355));
  nor2   g0291(.a(n352), .b(n355), .O(n356));
  nor2   g0292(.a(n356), .b(n354), .O(n357));
  inv1   g0293(.a(n357), .O(n358));
  nor2   g0294(.a(n358), .b(n303), .O(n359));
  inv1   g0295(.a(n303), .O(n360));
  nor2   g0296(.a(n357), .b(n360), .O(n361));
  nor2   g0297(.a(n361), .b(n359), .O(n362));
  inv1   g0298(.a(n362), .O(n363));
  nor2   g0299(.a(n363), .b(n302), .O(n364));
  inv1   g0300(.a(n302), .O(n365));
  nor2   g0301(.a(n362), .b(n365), .O(n366));
  nor2   g0302(.a(n366), .b(n364), .O(n367));
  inv1   g0303(.a(n367), .O(n368));
  nor2   g0304(.a(n368), .b(n301), .O(n369));
  inv1   g0305(.a(n301), .O(n370));
  nor2   g0306(.a(n367), .b(n370), .O(n371));
  nor2   g0307(.a(n371), .b(n369), .O(n372));
  inv1   g0308(.a(n372), .O(n373));
  nor2   g0309(.a(n373), .b(n300), .O(n374));
  inv1   g0310(.a(n300), .O(n375));
  nor2   g0311(.a(n372), .b(n375), .O(n376));
  nor2   g0312(.a(n376), .b(n374), .O(n377));
  inv1   g0313(.a(n377), .O(G3552gat));
  inv1   g0314(.a(G409gat), .O(n379));
  nor2   g0315(.a(n379), .b(n65), .O(n380));
  nor2   g0316(.a(n374), .b(n369), .O(n381));
  nor2   g0317(.a(n299), .b(n68), .O(n382));
  nor2   g0318(.a(n364), .b(n359), .O(n383));
  nor2   g0319(.a(n231), .b(n82), .O(n384));
  nor2   g0320(.a(n354), .b(n349), .O(n385));
  nor2   g0321(.a(n175), .b(n104), .O(n386));
  nor2   g0322(.a(n344), .b(n339), .O(n387));
  nor2   g0323(.a(n131), .b(n138), .O(n388));
  nor2   g0324(.a(n334), .b(n329), .O(n389));
  nor2   g0325(.a(n100), .b(n184), .O(n390));
  nor2   g0326(.a(n319), .b(n318), .O(n391));
  nor2   g0327(.a(n391), .b(n323), .O(n392));
  nor2   g0328(.a(n78), .b(n242), .O(n393));
  inv1   g0329(.a(G137gat), .O(n394));
  nor2   g0330(.a(n66), .b(n394), .O(n395));
  inv1   g0331(.a(n395), .O(n396));
  nor2   g0332(.a(n71), .b(n312), .O(n397));
  inv1   g0333(.a(n397), .O(n398));
  nor2   g0334(.a(n398), .b(G103gat), .O(n399));
  nor2   g0335(.a(n399), .b(n396), .O(n400));
  nor2   g0336(.a(n398), .b(n395), .O(n401));
  inv1   g0337(.a(n401), .O(n402));
  nor2   g0338(.a(n402), .b(n243), .O(n403));
  nor2   g0339(.a(n403), .b(n400), .O(n404));
  nor2   g0340(.a(n404), .b(n393), .O(n405));
  inv1   g0341(.a(n393), .O(n406));
  inv1   g0342(.a(n404), .O(n407));
  nor2   g0343(.a(n407), .b(n406), .O(n408));
  nor2   g0344(.a(n408), .b(n405), .O(n409));
  inv1   g0345(.a(n409), .O(n410));
  nor2   g0346(.a(n410), .b(n392), .O(n411));
  inv1   g0347(.a(n392), .O(n412));
  nor2   g0348(.a(n409), .b(n412), .O(n413));
  nor2   g0349(.a(n413), .b(n411), .O(n414));
  inv1   g0350(.a(n414), .O(n415));
  nor2   g0351(.a(n415), .b(n390), .O(n416));
  inv1   g0352(.a(n390), .O(n417));
  nor2   g0353(.a(n414), .b(n417), .O(n418));
  nor2   g0354(.a(n418), .b(n416), .O(n419));
  inv1   g0355(.a(n419), .O(n420));
  nor2   g0356(.a(n420), .b(n389), .O(n421));
  inv1   g0357(.a(n389), .O(n422));
  nor2   g0358(.a(n419), .b(n422), .O(n423));
  nor2   g0359(.a(n423), .b(n421), .O(n424));
  inv1   g0360(.a(n424), .O(n425));
  nor2   g0361(.a(n425), .b(n388), .O(n426));
  inv1   g0362(.a(n388), .O(n427));
  nor2   g0363(.a(n424), .b(n427), .O(n428));
  nor2   g0364(.a(n428), .b(n426), .O(n429));
  inv1   g0365(.a(n429), .O(n430));
  nor2   g0366(.a(n430), .b(n387), .O(n431));
  inv1   g0367(.a(n387), .O(n432));
  nor2   g0368(.a(n429), .b(n432), .O(n433));
  nor2   g0369(.a(n433), .b(n431), .O(n434));
  inv1   g0370(.a(n434), .O(n435));
  nor2   g0371(.a(n435), .b(n386), .O(n436));
  inv1   g0372(.a(n386), .O(n437));
  nor2   g0373(.a(n434), .b(n437), .O(n438));
  nor2   g0374(.a(n438), .b(n436), .O(n439));
  inv1   g0375(.a(n439), .O(n440));
  nor2   g0376(.a(n440), .b(n385), .O(n441));
  inv1   g0377(.a(n385), .O(n442));
  nor2   g0378(.a(n439), .b(n442), .O(n443));
  nor2   g0379(.a(n443), .b(n441), .O(n444));
  inv1   g0380(.a(n444), .O(n445));
  nor2   g0381(.a(n445), .b(n384), .O(n446));
  inv1   g0382(.a(n384), .O(n447));
  nor2   g0383(.a(n444), .b(n447), .O(n448));
  nor2   g0384(.a(n448), .b(n446), .O(n449));
  inv1   g0385(.a(n449), .O(n450));
  nor2   g0386(.a(n450), .b(n383), .O(n451));
  inv1   g0387(.a(n383), .O(n452));
  nor2   g0388(.a(n449), .b(n452), .O(n453));
  nor2   g0389(.a(n453), .b(n451), .O(n454));
  inv1   g0390(.a(n454), .O(n455));
  nor2   g0391(.a(n455), .b(n382), .O(n456));
  inv1   g0392(.a(n382), .O(n457));
  nor2   g0393(.a(n454), .b(n457), .O(n458));
  nor2   g0394(.a(n458), .b(n456), .O(n459));
  inv1   g0395(.a(n459), .O(n460));
  nor2   g0396(.a(n460), .b(n381), .O(n461));
  inv1   g0397(.a(n381), .O(n462));
  nor2   g0398(.a(n459), .b(n462), .O(n463));
  nor2   g0399(.a(n463), .b(n461), .O(n464));
  inv1   g0400(.a(n464), .O(n465));
  nor2   g0401(.a(n465), .b(n380), .O(n466));
  inv1   g0402(.a(n380), .O(n467));
  nor2   g0403(.a(n464), .b(n467), .O(n468));
  nor2   g0404(.a(n468), .b(n466), .O(n469));
  inv1   g0405(.a(n469), .O(G3895gat));
  inv1   g0406(.a(G426gat), .O(n471));
  nor2   g0407(.a(n471), .b(n65), .O(n472));
  nor2   g0408(.a(n466), .b(n461), .O(n473));
  nor2   g0409(.a(n379), .b(n68), .O(n474));
  nor2   g0410(.a(n456), .b(n451), .O(n475));
  nor2   g0411(.a(n299), .b(n82), .O(n476));
  nor2   g0412(.a(n446), .b(n441), .O(n477));
  nor2   g0413(.a(n231), .b(n104), .O(n478));
  nor2   g0414(.a(n436), .b(n431), .O(n479));
  nor2   g0415(.a(n175), .b(n138), .O(n480));
  nor2   g0416(.a(n426), .b(n421), .O(n481));
  nor2   g0417(.a(n131), .b(n184), .O(n482));
  nor2   g0418(.a(n416), .b(n411), .O(n483));
  nor2   g0419(.a(n100), .b(n242), .O(n484));
  nor2   g0420(.a(n401), .b(n400), .O(n485));
  nor2   g0421(.a(n485), .b(n405), .O(n486));
  nor2   g0422(.a(n78), .b(n312), .O(n487));
  inv1   g0423(.a(G154gat), .O(n488));
  nor2   g0424(.a(n66), .b(n488), .O(n489));
  inv1   g0425(.a(n489), .O(n490));
  nor2   g0426(.a(n71), .b(n394), .O(n491));
  inv1   g0427(.a(n491), .O(n492));
  nor2   g0428(.a(n492), .b(G120gat), .O(n493));
  nor2   g0429(.a(n493), .b(n490), .O(n494));
  nor2   g0430(.a(n492), .b(n489), .O(n495));
  inv1   g0431(.a(n495), .O(n496));
  nor2   g0432(.a(n496), .b(n313), .O(n497));
  nor2   g0433(.a(n497), .b(n494), .O(n498));
  nor2   g0434(.a(n498), .b(n487), .O(n499));
  inv1   g0435(.a(n487), .O(n500));
  inv1   g0436(.a(n498), .O(n501));
  nor2   g0437(.a(n501), .b(n500), .O(n502));
  nor2   g0438(.a(n502), .b(n499), .O(n503));
  inv1   g0439(.a(n503), .O(n504));
  nor2   g0440(.a(n504), .b(n486), .O(n505));
  inv1   g0441(.a(n486), .O(n506));
  nor2   g0442(.a(n503), .b(n506), .O(n507));
  nor2   g0443(.a(n507), .b(n505), .O(n508));
  inv1   g0444(.a(n508), .O(n509));
  nor2   g0445(.a(n509), .b(n484), .O(n510));
  inv1   g0446(.a(n484), .O(n511));
  nor2   g0447(.a(n508), .b(n511), .O(n512));
  nor2   g0448(.a(n512), .b(n510), .O(n513));
  inv1   g0449(.a(n513), .O(n514));
  nor2   g0450(.a(n514), .b(n483), .O(n515));
  inv1   g0451(.a(n483), .O(n516));
  nor2   g0452(.a(n513), .b(n516), .O(n517));
  nor2   g0453(.a(n517), .b(n515), .O(n518));
  inv1   g0454(.a(n518), .O(n519));
  nor2   g0455(.a(n519), .b(n482), .O(n520));
  inv1   g0456(.a(n482), .O(n521));
  nor2   g0457(.a(n518), .b(n521), .O(n522));
  nor2   g0458(.a(n522), .b(n520), .O(n523));
  inv1   g0459(.a(n523), .O(n524));
  nor2   g0460(.a(n524), .b(n481), .O(n525));
  inv1   g0461(.a(n481), .O(n526));
  nor2   g0462(.a(n523), .b(n526), .O(n527));
  nor2   g0463(.a(n527), .b(n525), .O(n528));
  inv1   g0464(.a(n528), .O(n529));
  nor2   g0465(.a(n529), .b(n480), .O(n530));
  inv1   g0466(.a(n480), .O(n531));
  nor2   g0467(.a(n528), .b(n531), .O(n532));
  nor2   g0468(.a(n532), .b(n530), .O(n533));
  inv1   g0469(.a(n533), .O(n534));
  nor2   g0470(.a(n534), .b(n479), .O(n535));
  inv1   g0471(.a(n479), .O(n536));
  nor2   g0472(.a(n533), .b(n536), .O(n537));
  nor2   g0473(.a(n537), .b(n535), .O(n538));
  inv1   g0474(.a(n538), .O(n539));
  nor2   g0475(.a(n539), .b(n478), .O(n540));
  inv1   g0476(.a(n478), .O(n541));
  nor2   g0477(.a(n538), .b(n541), .O(n542));
  nor2   g0478(.a(n542), .b(n540), .O(n543));
  inv1   g0479(.a(n543), .O(n544));
  nor2   g0480(.a(n544), .b(n477), .O(n545));
  inv1   g0481(.a(n477), .O(n546));
  nor2   g0482(.a(n543), .b(n546), .O(n547));
  nor2   g0483(.a(n547), .b(n545), .O(n548));
  inv1   g0484(.a(n548), .O(n549));
  nor2   g0485(.a(n549), .b(n476), .O(n550));
  inv1   g0486(.a(n476), .O(n551));
  nor2   g0487(.a(n548), .b(n551), .O(n552));
  nor2   g0488(.a(n552), .b(n550), .O(n553));
  inv1   g0489(.a(n553), .O(n554));
  nor2   g0490(.a(n554), .b(n475), .O(n555));
  inv1   g0491(.a(n475), .O(n556));
  nor2   g0492(.a(n553), .b(n556), .O(n557));
  nor2   g0493(.a(n557), .b(n555), .O(n558));
  inv1   g0494(.a(n558), .O(n559));
  nor2   g0495(.a(n559), .b(n474), .O(n560));
  inv1   g0496(.a(n474), .O(n561));
  nor2   g0497(.a(n558), .b(n561), .O(n562));
  nor2   g0498(.a(n562), .b(n560), .O(n563));
  inv1   g0499(.a(n563), .O(n564));
  nor2   g0500(.a(n564), .b(n473), .O(n565));
  inv1   g0501(.a(n473), .O(n566));
  nor2   g0502(.a(n563), .b(n566), .O(n567));
  nor2   g0503(.a(n567), .b(n565), .O(n568));
  inv1   g0504(.a(n568), .O(n569));
  nor2   g0505(.a(n569), .b(n472), .O(n570));
  inv1   g0506(.a(n472), .O(n571));
  nor2   g0507(.a(n568), .b(n571), .O(n572));
  nor2   g0508(.a(n572), .b(n570), .O(n573));
  inv1   g0509(.a(n573), .O(G4241gat));
  inv1   g0510(.a(G443gat), .O(n575));
  nor2   g0511(.a(n575), .b(n65), .O(n576));
  nor2   g0512(.a(n570), .b(n565), .O(n577));
  nor2   g0513(.a(n471), .b(n68), .O(n578));
  nor2   g0514(.a(n560), .b(n555), .O(n579));
  nor2   g0515(.a(n379), .b(n82), .O(n580));
  nor2   g0516(.a(n550), .b(n545), .O(n581));
  nor2   g0517(.a(n299), .b(n104), .O(n582));
  nor2   g0518(.a(n540), .b(n535), .O(n583));
  nor2   g0519(.a(n231), .b(n138), .O(n584));
  nor2   g0520(.a(n530), .b(n525), .O(n585));
  nor2   g0521(.a(n175), .b(n184), .O(n586));
  nor2   g0522(.a(n520), .b(n515), .O(n587));
  nor2   g0523(.a(n131), .b(n242), .O(n588));
  nor2   g0524(.a(n510), .b(n505), .O(n589));
  nor2   g0525(.a(n100), .b(n312), .O(n590));
  nor2   g0526(.a(n495), .b(n494), .O(n591));
  nor2   g0527(.a(n591), .b(n499), .O(n592));
  nor2   g0528(.a(n78), .b(n394), .O(n593));
  inv1   g0529(.a(G171gat), .O(n594));
  nor2   g0530(.a(n66), .b(n594), .O(n595));
  inv1   g0531(.a(n595), .O(n596));
  nor2   g0532(.a(n71), .b(n488), .O(n597));
  inv1   g0533(.a(n597), .O(n598));
  nor2   g0534(.a(n598), .b(G137gat), .O(n599));
  nor2   g0535(.a(n599), .b(n596), .O(n600));
  nor2   g0536(.a(n598), .b(n595), .O(n601));
  inv1   g0537(.a(n601), .O(n602));
  nor2   g0538(.a(n602), .b(n395), .O(n603));
  nor2   g0539(.a(n603), .b(n600), .O(n604));
  nor2   g0540(.a(n604), .b(n593), .O(n605));
  inv1   g0541(.a(n593), .O(n606));
  inv1   g0542(.a(n604), .O(n607));
  nor2   g0543(.a(n607), .b(n606), .O(n608));
  nor2   g0544(.a(n608), .b(n605), .O(n609));
  inv1   g0545(.a(n609), .O(n610));
  nor2   g0546(.a(n610), .b(n592), .O(n611));
  inv1   g0547(.a(n592), .O(n612));
  nor2   g0548(.a(n609), .b(n612), .O(n613));
  nor2   g0549(.a(n613), .b(n611), .O(n614));
  inv1   g0550(.a(n614), .O(n615));
  nor2   g0551(.a(n615), .b(n590), .O(n616));
  inv1   g0552(.a(n590), .O(n617));
  nor2   g0553(.a(n614), .b(n617), .O(n618));
  nor2   g0554(.a(n618), .b(n616), .O(n619));
  inv1   g0555(.a(n619), .O(n620));
  nor2   g0556(.a(n620), .b(n589), .O(n621));
  inv1   g0557(.a(n589), .O(n622));
  nor2   g0558(.a(n619), .b(n622), .O(n623));
  nor2   g0559(.a(n623), .b(n621), .O(n624));
  inv1   g0560(.a(n624), .O(n625));
  nor2   g0561(.a(n625), .b(n588), .O(n626));
  inv1   g0562(.a(n588), .O(n627));
  nor2   g0563(.a(n624), .b(n627), .O(n628));
  nor2   g0564(.a(n628), .b(n626), .O(n629));
  inv1   g0565(.a(n629), .O(n630));
  nor2   g0566(.a(n630), .b(n587), .O(n631));
  inv1   g0567(.a(n587), .O(n632));
  nor2   g0568(.a(n629), .b(n632), .O(n633));
  nor2   g0569(.a(n633), .b(n631), .O(n634));
  inv1   g0570(.a(n634), .O(n635));
  nor2   g0571(.a(n635), .b(n586), .O(n636));
  inv1   g0572(.a(n586), .O(n637));
  nor2   g0573(.a(n634), .b(n637), .O(n638));
  nor2   g0574(.a(n638), .b(n636), .O(n639));
  inv1   g0575(.a(n639), .O(n640));
  nor2   g0576(.a(n640), .b(n585), .O(n641));
  inv1   g0577(.a(n585), .O(n642));
  nor2   g0578(.a(n639), .b(n642), .O(n643));
  nor2   g0579(.a(n643), .b(n641), .O(n644));
  inv1   g0580(.a(n644), .O(n645));
  nor2   g0581(.a(n645), .b(n584), .O(n646));
  inv1   g0582(.a(n584), .O(n647));
  nor2   g0583(.a(n644), .b(n647), .O(n648));
  nor2   g0584(.a(n648), .b(n646), .O(n649));
  inv1   g0585(.a(n649), .O(n650));
  nor2   g0586(.a(n650), .b(n583), .O(n651));
  inv1   g0587(.a(n583), .O(n652));
  nor2   g0588(.a(n649), .b(n652), .O(n653));
  nor2   g0589(.a(n653), .b(n651), .O(n654));
  inv1   g0590(.a(n654), .O(n655));
  nor2   g0591(.a(n655), .b(n582), .O(n656));
  inv1   g0592(.a(n582), .O(n657));
  nor2   g0593(.a(n654), .b(n657), .O(n658));
  nor2   g0594(.a(n658), .b(n656), .O(n659));
  inv1   g0595(.a(n659), .O(n660));
  nor2   g0596(.a(n660), .b(n581), .O(n661));
  inv1   g0597(.a(n581), .O(n662));
  nor2   g0598(.a(n659), .b(n662), .O(n663));
  nor2   g0599(.a(n663), .b(n661), .O(n664));
  inv1   g0600(.a(n664), .O(n665));
  nor2   g0601(.a(n665), .b(n580), .O(n666));
  inv1   g0602(.a(n580), .O(n667));
  nor2   g0603(.a(n664), .b(n667), .O(n668));
  nor2   g0604(.a(n668), .b(n666), .O(n669));
  inv1   g0605(.a(n669), .O(n670));
  nor2   g0606(.a(n670), .b(n579), .O(n671));
  inv1   g0607(.a(n579), .O(n672));
  nor2   g0608(.a(n669), .b(n672), .O(n673));
  nor2   g0609(.a(n673), .b(n671), .O(n674));
  inv1   g0610(.a(n674), .O(n675));
  nor2   g0611(.a(n675), .b(n578), .O(n676));
  inv1   g0612(.a(n578), .O(n677));
  nor2   g0613(.a(n674), .b(n677), .O(n678));
  nor2   g0614(.a(n678), .b(n676), .O(n679));
  inv1   g0615(.a(n679), .O(n680));
  nor2   g0616(.a(n680), .b(n577), .O(n681));
  inv1   g0617(.a(n577), .O(n682));
  nor2   g0618(.a(n679), .b(n682), .O(n683));
  nor2   g0619(.a(n683), .b(n681), .O(n684));
  inv1   g0620(.a(n684), .O(n685));
  nor2   g0621(.a(n685), .b(n576), .O(n686));
  inv1   g0622(.a(n576), .O(n687));
  nor2   g0623(.a(n684), .b(n687), .O(n688));
  nor2   g0624(.a(n688), .b(n686), .O(n689));
  inv1   g0625(.a(n689), .O(G4591gat));
  inv1   g0626(.a(G460gat), .O(n691));
  nor2   g0627(.a(n691), .b(n65), .O(n692));
  nor2   g0628(.a(n686), .b(n681), .O(n693));
  nor2   g0629(.a(n575), .b(n68), .O(n694));
  nor2   g0630(.a(n676), .b(n671), .O(n695));
  nor2   g0631(.a(n471), .b(n82), .O(n696));
  nor2   g0632(.a(n666), .b(n661), .O(n697));
  nor2   g0633(.a(n379), .b(n104), .O(n698));
  nor2   g0634(.a(n656), .b(n651), .O(n699));
  nor2   g0635(.a(n299), .b(n138), .O(n700));
  nor2   g0636(.a(n646), .b(n641), .O(n701));
  nor2   g0637(.a(n231), .b(n184), .O(n702));
  nor2   g0638(.a(n636), .b(n631), .O(n703));
  nor2   g0639(.a(n175), .b(n242), .O(n704));
  nor2   g0640(.a(n626), .b(n621), .O(n705));
  nor2   g0641(.a(n131), .b(n312), .O(n706));
  nor2   g0642(.a(n616), .b(n611), .O(n707));
  nor2   g0643(.a(n100), .b(n394), .O(n708));
  nor2   g0644(.a(n601), .b(n600), .O(n709));
  nor2   g0645(.a(n709), .b(n605), .O(n710));
  nor2   g0646(.a(n78), .b(n488), .O(n711));
  inv1   g0647(.a(G188gat), .O(n712));
  nor2   g0648(.a(n66), .b(n712), .O(n713));
  inv1   g0649(.a(n713), .O(n714));
  nor2   g0650(.a(n71), .b(n594), .O(n715));
  inv1   g0651(.a(n715), .O(n716));
  nor2   g0652(.a(n716), .b(G154gat), .O(n717));
  nor2   g0653(.a(n717), .b(n714), .O(n718));
  nor2   g0654(.a(n716), .b(n713), .O(n719));
  inv1   g0655(.a(n719), .O(n720));
  nor2   g0656(.a(n720), .b(n489), .O(n721));
  nor2   g0657(.a(n721), .b(n718), .O(n722));
  nor2   g0658(.a(n722), .b(n711), .O(n723));
  inv1   g0659(.a(n711), .O(n724));
  inv1   g0660(.a(n722), .O(n725));
  nor2   g0661(.a(n725), .b(n724), .O(n726));
  nor2   g0662(.a(n726), .b(n723), .O(n727));
  inv1   g0663(.a(n727), .O(n728));
  nor2   g0664(.a(n728), .b(n710), .O(n729));
  inv1   g0665(.a(n710), .O(n730));
  nor2   g0666(.a(n727), .b(n730), .O(n731));
  nor2   g0667(.a(n731), .b(n729), .O(n732));
  inv1   g0668(.a(n732), .O(n733));
  nor2   g0669(.a(n733), .b(n708), .O(n734));
  inv1   g0670(.a(n708), .O(n735));
  nor2   g0671(.a(n732), .b(n735), .O(n736));
  nor2   g0672(.a(n736), .b(n734), .O(n737));
  inv1   g0673(.a(n737), .O(n738));
  nor2   g0674(.a(n738), .b(n707), .O(n739));
  inv1   g0675(.a(n707), .O(n740));
  nor2   g0676(.a(n737), .b(n740), .O(n741));
  nor2   g0677(.a(n741), .b(n739), .O(n742));
  inv1   g0678(.a(n742), .O(n743));
  nor2   g0679(.a(n743), .b(n706), .O(n744));
  inv1   g0680(.a(n706), .O(n745));
  nor2   g0681(.a(n742), .b(n745), .O(n746));
  nor2   g0682(.a(n746), .b(n744), .O(n747));
  inv1   g0683(.a(n747), .O(n748));
  nor2   g0684(.a(n748), .b(n705), .O(n749));
  inv1   g0685(.a(n705), .O(n750));
  nor2   g0686(.a(n747), .b(n750), .O(n751));
  nor2   g0687(.a(n751), .b(n749), .O(n752));
  inv1   g0688(.a(n752), .O(n753));
  nor2   g0689(.a(n753), .b(n704), .O(n754));
  inv1   g0690(.a(n704), .O(n755));
  nor2   g0691(.a(n752), .b(n755), .O(n756));
  nor2   g0692(.a(n756), .b(n754), .O(n757));
  inv1   g0693(.a(n757), .O(n758));
  nor2   g0694(.a(n758), .b(n703), .O(n759));
  inv1   g0695(.a(n703), .O(n760));
  nor2   g0696(.a(n757), .b(n760), .O(n761));
  nor2   g0697(.a(n761), .b(n759), .O(n762));
  inv1   g0698(.a(n762), .O(n763));
  nor2   g0699(.a(n763), .b(n702), .O(n764));
  inv1   g0700(.a(n702), .O(n765));
  nor2   g0701(.a(n762), .b(n765), .O(n766));
  nor2   g0702(.a(n766), .b(n764), .O(n767));
  inv1   g0703(.a(n767), .O(n768));
  nor2   g0704(.a(n768), .b(n701), .O(n769));
  inv1   g0705(.a(n701), .O(n770));
  nor2   g0706(.a(n767), .b(n770), .O(n771));
  nor2   g0707(.a(n771), .b(n769), .O(n772));
  inv1   g0708(.a(n772), .O(n773));
  nor2   g0709(.a(n773), .b(n700), .O(n774));
  inv1   g0710(.a(n700), .O(n775));
  nor2   g0711(.a(n772), .b(n775), .O(n776));
  nor2   g0712(.a(n776), .b(n774), .O(n777));
  inv1   g0713(.a(n777), .O(n778));
  nor2   g0714(.a(n778), .b(n699), .O(n779));
  inv1   g0715(.a(n699), .O(n780));
  nor2   g0716(.a(n777), .b(n780), .O(n781));
  nor2   g0717(.a(n781), .b(n779), .O(n782));
  inv1   g0718(.a(n782), .O(n783));
  nor2   g0719(.a(n783), .b(n698), .O(n784));
  inv1   g0720(.a(n698), .O(n785));
  nor2   g0721(.a(n782), .b(n785), .O(n786));
  nor2   g0722(.a(n786), .b(n784), .O(n787));
  inv1   g0723(.a(n787), .O(n788));
  nor2   g0724(.a(n788), .b(n697), .O(n789));
  inv1   g0725(.a(n697), .O(n790));
  nor2   g0726(.a(n787), .b(n790), .O(n791));
  nor2   g0727(.a(n791), .b(n789), .O(n792));
  inv1   g0728(.a(n792), .O(n793));
  nor2   g0729(.a(n793), .b(n696), .O(n794));
  inv1   g0730(.a(n696), .O(n795));
  nor2   g0731(.a(n792), .b(n795), .O(n796));
  nor2   g0732(.a(n796), .b(n794), .O(n797));
  inv1   g0733(.a(n797), .O(n798));
  nor2   g0734(.a(n798), .b(n695), .O(n799));
  inv1   g0735(.a(n695), .O(n800));
  nor2   g0736(.a(n797), .b(n800), .O(n801));
  nor2   g0737(.a(n801), .b(n799), .O(n802));
  inv1   g0738(.a(n802), .O(n803));
  nor2   g0739(.a(n803), .b(n694), .O(n804));
  inv1   g0740(.a(n694), .O(n805));
  nor2   g0741(.a(n802), .b(n805), .O(n806));
  nor2   g0742(.a(n806), .b(n804), .O(n807));
  inv1   g0743(.a(n807), .O(n808));
  nor2   g0744(.a(n808), .b(n693), .O(n809));
  inv1   g0745(.a(n693), .O(n810));
  nor2   g0746(.a(n807), .b(n810), .O(n811));
  nor2   g0747(.a(n811), .b(n809), .O(n812));
  inv1   g0748(.a(n812), .O(n813));
  nor2   g0749(.a(n813), .b(n692), .O(n814));
  inv1   g0750(.a(n692), .O(n815));
  nor2   g0751(.a(n812), .b(n815), .O(n816));
  nor2   g0752(.a(n816), .b(n814), .O(n817));
  inv1   g0753(.a(n817), .O(G4946gat));
  inv1   g0754(.a(G477gat), .O(n819));
  nor2   g0755(.a(n819), .b(n65), .O(n820));
  nor2   g0756(.a(n814), .b(n809), .O(n821));
  nor2   g0757(.a(n691), .b(n68), .O(n822));
  nor2   g0758(.a(n804), .b(n799), .O(n823));
  nor2   g0759(.a(n575), .b(n82), .O(n824));
  nor2   g0760(.a(n794), .b(n789), .O(n825));
  nor2   g0761(.a(n471), .b(n104), .O(n826));
  nor2   g0762(.a(n784), .b(n779), .O(n827));
  nor2   g0763(.a(n379), .b(n138), .O(n828));
  nor2   g0764(.a(n774), .b(n769), .O(n829));
  nor2   g0765(.a(n299), .b(n184), .O(n830));
  nor2   g0766(.a(n764), .b(n759), .O(n831));
  nor2   g0767(.a(n231), .b(n242), .O(n832));
  nor2   g0768(.a(n754), .b(n749), .O(n833));
  nor2   g0769(.a(n175), .b(n312), .O(n834));
  nor2   g0770(.a(n744), .b(n739), .O(n835));
  nor2   g0771(.a(n131), .b(n394), .O(n836));
  nor2   g0772(.a(n734), .b(n729), .O(n837));
  nor2   g0773(.a(n100), .b(n488), .O(n838));
  nor2   g0774(.a(n719), .b(n718), .O(n839));
  nor2   g0775(.a(n839), .b(n723), .O(n840));
  nor2   g0776(.a(n78), .b(n594), .O(n841));
  inv1   g0777(.a(G205gat), .O(n842));
  nor2   g0778(.a(n66), .b(n842), .O(n843));
  inv1   g0779(.a(n843), .O(n844));
  nor2   g0780(.a(n71), .b(n712), .O(n845));
  inv1   g0781(.a(n845), .O(n846));
  nor2   g0782(.a(n846), .b(G171gat), .O(n847));
  nor2   g0783(.a(n847), .b(n844), .O(n848));
  nor2   g0784(.a(n846), .b(n843), .O(n849));
  inv1   g0785(.a(n849), .O(n850));
  nor2   g0786(.a(n850), .b(n595), .O(n851));
  nor2   g0787(.a(n851), .b(n848), .O(n852));
  nor2   g0788(.a(n852), .b(n841), .O(n853));
  inv1   g0789(.a(n841), .O(n854));
  inv1   g0790(.a(n852), .O(n855));
  nor2   g0791(.a(n855), .b(n854), .O(n856));
  nor2   g0792(.a(n856), .b(n853), .O(n857));
  inv1   g0793(.a(n857), .O(n858));
  nor2   g0794(.a(n858), .b(n840), .O(n859));
  inv1   g0795(.a(n840), .O(n860));
  nor2   g0796(.a(n857), .b(n860), .O(n861));
  nor2   g0797(.a(n861), .b(n859), .O(n862));
  inv1   g0798(.a(n862), .O(n863));
  nor2   g0799(.a(n863), .b(n838), .O(n864));
  inv1   g0800(.a(n838), .O(n865));
  nor2   g0801(.a(n862), .b(n865), .O(n866));
  nor2   g0802(.a(n866), .b(n864), .O(n867));
  inv1   g0803(.a(n867), .O(n868));
  nor2   g0804(.a(n868), .b(n837), .O(n869));
  inv1   g0805(.a(n837), .O(n870));
  nor2   g0806(.a(n867), .b(n870), .O(n871));
  nor2   g0807(.a(n871), .b(n869), .O(n872));
  inv1   g0808(.a(n872), .O(n873));
  nor2   g0809(.a(n873), .b(n836), .O(n874));
  inv1   g0810(.a(n836), .O(n875));
  nor2   g0811(.a(n872), .b(n875), .O(n876));
  nor2   g0812(.a(n876), .b(n874), .O(n877));
  inv1   g0813(.a(n877), .O(n878));
  nor2   g0814(.a(n878), .b(n835), .O(n879));
  inv1   g0815(.a(n835), .O(n880));
  nor2   g0816(.a(n877), .b(n880), .O(n881));
  nor2   g0817(.a(n881), .b(n879), .O(n882));
  inv1   g0818(.a(n882), .O(n883));
  nor2   g0819(.a(n883), .b(n834), .O(n884));
  inv1   g0820(.a(n834), .O(n885));
  nor2   g0821(.a(n882), .b(n885), .O(n886));
  nor2   g0822(.a(n886), .b(n884), .O(n887));
  inv1   g0823(.a(n887), .O(n888));
  nor2   g0824(.a(n888), .b(n833), .O(n889));
  inv1   g0825(.a(n833), .O(n890));
  nor2   g0826(.a(n887), .b(n890), .O(n891));
  nor2   g0827(.a(n891), .b(n889), .O(n892));
  inv1   g0828(.a(n892), .O(n893));
  nor2   g0829(.a(n893), .b(n832), .O(n894));
  inv1   g0830(.a(n832), .O(n895));
  nor2   g0831(.a(n892), .b(n895), .O(n896));
  nor2   g0832(.a(n896), .b(n894), .O(n897));
  inv1   g0833(.a(n897), .O(n898));
  nor2   g0834(.a(n898), .b(n831), .O(n899));
  inv1   g0835(.a(n831), .O(n900));
  nor2   g0836(.a(n897), .b(n900), .O(n901));
  nor2   g0837(.a(n901), .b(n899), .O(n902));
  inv1   g0838(.a(n902), .O(n903));
  nor2   g0839(.a(n903), .b(n830), .O(n904));
  inv1   g0840(.a(n830), .O(n905));
  nor2   g0841(.a(n902), .b(n905), .O(n906));
  nor2   g0842(.a(n906), .b(n904), .O(n907));
  inv1   g0843(.a(n907), .O(n908));
  nor2   g0844(.a(n908), .b(n829), .O(n909));
  inv1   g0845(.a(n829), .O(n910));
  nor2   g0846(.a(n907), .b(n910), .O(n911));
  nor2   g0847(.a(n911), .b(n909), .O(n912));
  inv1   g0848(.a(n912), .O(n913));
  nor2   g0849(.a(n913), .b(n828), .O(n914));
  inv1   g0850(.a(n828), .O(n915));
  nor2   g0851(.a(n912), .b(n915), .O(n916));
  nor2   g0852(.a(n916), .b(n914), .O(n917));
  inv1   g0853(.a(n917), .O(n918));
  nor2   g0854(.a(n918), .b(n827), .O(n919));
  inv1   g0855(.a(n827), .O(n920));
  nor2   g0856(.a(n917), .b(n920), .O(n921));
  nor2   g0857(.a(n921), .b(n919), .O(n922));
  inv1   g0858(.a(n922), .O(n923));
  nor2   g0859(.a(n923), .b(n826), .O(n924));
  inv1   g0860(.a(n826), .O(n925));
  nor2   g0861(.a(n922), .b(n925), .O(n926));
  nor2   g0862(.a(n926), .b(n924), .O(n927));
  inv1   g0863(.a(n927), .O(n928));
  nor2   g0864(.a(n928), .b(n825), .O(n929));
  inv1   g0865(.a(n825), .O(n930));
  nor2   g0866(.a(n927), .b(n930), .O(n931));
  nor2   g0867(.a(n931), .b(n929), .O(n932));
  inv1   g0868(.a(n932), .O(n933));
  nor2   g0869(.a(n933), .b(n824), .O(n934));
  inv1   g0870(.a(n824), .O(n935));
  nor2   g0871(.a(n932), .b(n935), .O(n936));
  nor2   g0872(.a(n936), .b(n934), .O(n937));
  inv1   g0873(.a(n937), .O(n938));
  nor2   g0874(.a(n938), .b(n823), .O(n939));
  inv1   g0875(.a(n823), .O(n940));
  nor2   g0876(.a(n937), .b(n940), .O(n941));
  nor2   g0877(.a(n941), .b(n939), .O(n942));
  inv1   g0878(.a(n942), .O(n943));
  nor2   g0879(.a(n943), .b(n822), .O(n944));
  inv1   g0880(.a(n822), .O(n945));
  nor2   g0881(.a(n942), .b(n945), .O(n946));
  nor2   g0882(.a(n946), .b(n944), .O(n947));
  inv1   g0883(.a(n947), .O(n948));
  nor2   g0884(.a(n948), .b(n821), .O(n949));
  inv1   g0885(.a(n821), .O(n950));
  nor2   g0886(.a(n947), .b(n950), .O(n951));
  nor2   g0887(.a(n951), .b(n949), .O(n952));
  inv1   g0888(.a(n952), .O(n953));
  nor2   g0889(.a(n953), .b(n820), .O(n954));
  inv1   g0890(.a(n820), .O(n955));
  nor2   g0891(.a(n952), .b(n955), .O(n956));
  nor2   g0892(.a(n956), .b(n954), .O(n957));
  inv1   g0893(.a(n957), .O(G5308gat));
  inv1   g0894(.a(G494gat), .O(n959));
  nor2   g0895(.a(n959), .b(n65), .O(n960));
  nor2   g0896(.a(n954), .b(n949), .O(n961));
  nor2   g0897(.a(n819), .b(n68), .O(n962));
  nor2   g0898(.a(n944), .b(n939), .O(n963));
  nor2   g0899(.a(n691), .b(n82), .O(n964));
  nor2   g0900(.a(n934), .b(n929), .O(n965));
  nor2   g0901(.a(n575), .b(n104), .O(n966));
  nor2   g0902(.a(n924), .b(n919), .O(n967));
  nor2   g0903(.a(n471), .b(n138), .O(n968));
  nor2   g0904(.a(n914), .b(n909), .O(n969));
  nor2   g0905(.a(n379), .b(n184), .O(n970));
  nor2   g0906(.a(n904), .b(n899), .O(n971));
  nor2   g0907(.a(n299), .b(n242), .O(n972));
  nor2   g0908(.a(n894), .b(n889), .O(n973));
  nor2   g0909(.a(n231), .b(n312), .O(n974));
  nor2   g0910(.a(n884), .b(n879), .O(n975));
  nor2   g0911(.a(n175), .b(n394), .O(n976));
  nor2   g0912(.a(n874), .b(n869), .O(n977));
  nor2   g0913(.a(n131), .b(n488), .O(n978));
  nor2   g0914(.a(n864), .b(n859), .O(n979));
  nor2   g0915(.a(n100), .b(n594), .O(n980));
  nor2   g0916(.a(n849), .b(n848), .O(n981));
  nor2   g0917(.a(n981), .b(n853), .O(n982));
  nor2   g0918(.a(n78), .b(n712), .O(n983));
  inv1   g0919(.a(G222gat), .O(n984));
  nor2   g0920(.a(n66), .b(n984), .O(n985));
  inv1   g0921(.a(n985), .O(n986));
  nor2   g0922(.a(n71), .b(n842), .O(n987));
  inv1   g0923(.a(n987), .O(n988));
  nor2   g0924(.a(n988), .b(G188gat), .O(n989));
  nor2   g0925(.a(n989), .b(n986), .O(n990));
  nor2   g0926(.a(n988), .b(n985), .O(n991));
  inv1   g0927(.a(n991), .O(n992));
  nor2   g0928(.a(n992), .b(n713), .O(n993));
  nor2   g0929(.a(n993), .b(n990), .O(n994));
  nor2   g0930(.a(n994), .b(n983), .O(n995));
  inv1   g0931(.a(n983), .O(n996));
  inv1   g0932(.a(n994), .O(n997));
  nor2   g0933(.a(n997), .b(n996), .O(n998));
  nor2   g0934(.a(n998), .b(n995), .O(n999));
  inv1   g0935(.a(n999), .O(n1000));
  nor2   g0936(.a(n1000), .b(n982), .O(n1001));
  inv1   g0937(.a(n982), .O(n1002));
  nor2   g0938(.a(n999), .b(n1002), .O(n1003));
  nor2   g0939(.a(n1003), .b(n1001), .O(n1004));
  inv1   g0940(.a(n1004), .O(n1005));
  nor2   g0941(.a(n1005), .b(n980), .O(n1006));
  inv1   g0942(.a(n980), .O(n1007));
  nor2   g0943(.a(n1004), .b(n1007), .O(n1008));
  nor2   g0944(.a(n1008), .b(n1006), .O(n1009));
  inv1   g0945(.a(n1009), .O(n1010));
  nor2   g0946(.a(n1010), .b(n979), .O(n1011));
  inv1   g0947(.a(n979), .O(n1012));
  nor2   g0948(.a(n1009), .b(n1012), .O(n1013));
  nor2   g0949(.a(n1013), .b(n1011), .O(n1014));
  inv1   g0950(.a(n1014), .O(n1015));
  nor2   g0951(.a(n1015), .b(n978), .O(n1016));
  inv1   g0952(.a(n978), .O(n1017));
  nor2   g0953(.a(n1014), .b(n1017), .O(n1018));
  nor2   g0954(.a(n1018), .b(n1016), .O(n1019));
  inv1   g0955(.a(n1019), .O(n1020));
  nor2   g0956(.a(n1020), .b(n977), .O(n1021));
  inv1   g0957(.a(n977), .O(n1022));
  nor2   g0958(.a(n1019), .b(n1022), .O(n1023));
  nor2   g0959(.a(n1023), .b(n1021), .O(n1024));
  inv1   g0960(.a(n1024), .O(n1025));
  nor2   g0961(.a(n1025), .b(n976), .O(n1026));
  inv1   g0962(.a(n976), .O(n1027));
  nor2   g0963(.a(n1024), .b(n1027), .O(n1028));
  nor2   g0964(.a(n1028), .b(n1026), .O(n1029));
  inv1   g0965(.a(n1029), .O(n1030));
  nor2   g0966(.a(n1030), .b(n975), .O(n1031));
  inv1   g0967(.a(n975), .O(n1032));
  nor2   g0968(.a(n1029), .b(n1032), .O(n1033));
  nor2   g0969(.a(n1033), .b(n1031), .O(n1034));
  inv1   g0970(.a(n1034), .O(n1035));
  nor2   g0971(.a(n1035), .b(n974), .O(n1036));
  inv1   g0972(.a(n974), .O(n1037));
  nor2   g0973(.a(n1034), .b(n1037), .O(n1038));
  nor2   g0974(.a(n1038), .b(n1036), .O(n1039));
  inv1   g0975(.a(n1039), .O(n1040));
  nor2   g0976(.a(n1040), .b(n973), .O(n1041));
  inv1   g0977(.a(n973), .O(n1042));
  nor2   g0978(.a(n1039), .b(n1042), .O(n1043));
  nor2   g0979(.a(n1043), .b(n1041), .O(n1044));
  inv1   g0980(.a(n1044), .O(n1045));
  nor2   g0981(.a(n1045), .b(n972), .O(n1046));
  inv1   g0982(.a(n972), .O(n1047));
  nor2   g0983(.a(n1044), .b(n1047), .O(n1048));
  nor2   g0984(.a(n1048), .b(n1046), .O(n1049));
  inv1   g0985(.a(n1049), .O(n1050));
  nor2   g0986(.a(n1050), .b(n971), .O(n1051));
  inv1   g0987(.a(n971), .O(n1052));
  nor2   g0988(.a(n1049), .b(n1052), .O(n1053));
  nor2   g0989(.a(n1053), .b(n1051), .O(n1054));
  inv1   g0990(.a(n1054), .O(n1055));
  nor2   g0991(.a(n1055), .b(n970), .O(n1056));
  inv1   g0992(.a(n970), .O(n1057));
  nor2   g0993(.a(n1054), .b(n1057), .O(n1058));
  nor2   g0994(.a(n1058), .b(n1056), .O(n1059));
  inv1   g0995(.a(n1059), .O(n1060));
  nor2   g0996(.a(n1060), .b(n969), .O(n1061));
  inv1   g0997(.a(n969), .O(n1062));
  nor2   g0998(.a(n1059), .b(n1062), .O(n1063));
  nor2   g0999(.a(n1063), .b(n1061), .O(n1064));
  inv1   g1000(.a(n1064), .O(n1065));
  nor2   g1001(.a(n1065), .b(n968), .O(n1066));
  inv1   g1002(.a(n968), .O(n1067));
  nor2   g1003(.a(n1064), .b(n1067), .O(n1068));
  nor2   g1004(.a(n1068), .b(n1066), .O(n1069));
  inv1   g1005(.a(n1069), .O(n1070));
  nor2   g1006(.a(n1070), .b(n967), .O(n1071));
  inv1   g1007(.a(n967), .O(n1072));
  nor2   g1008(.a(n1069), .b(n1072), .O(n1073));
  nor2   g1009(.a(n1073), .b(n1071), .O(n1074));
  inv1   g1010(.a(n1074), .O(n1075));
  nor2   g1011(.a(n1075), .b(n966), .O(n1076));
  inv1   g1012(.a(n966), .O(n1077));
  nor2   g1013(.a(n1074), .b(n1077), .O(n1078));
  nor2   g1014(.a(n1078), .b(n1076), .O(n1079));
  inv1   g1015(.a(n1079), .O(n1080));
  nor2   g1016(.a(n1080), .b(n965), .O(n1081));
  inv1   g1017(.a(n965), .O(n1082));
  nor2   g1018(.a(n1079), .b(n1082), .O(n1083));
  nor2   g1019(.a(n1083), .b(n1081), .O(n1084));
  inv1   g1020(.a(n1084), .O(n1085));
  nor2   g1021(.a(n1085), .b(n964), .O(n1086));
  inv1   g1022(.a(n964), .O(n1087));
  nor2   g1023(.a(n1084), .b(n1087), .O(n1088));
  nor2   g1024(.a(n1088), .b(n1086), .O(n1089));
  inv1   g1025(.a(n1089), .O(n1090));
  nor2   g1026(.a(n1090), .b(n963), .O(n1091));
  inv1   g1027(.a(n963), .O(n1092));
  nor2   g1028(.a(n1089), .b(n1092), .O(n1093));
  nor2   g1029(.a(n1093), .b(n1091), .O(n1094));
  inv1   g1030(.a(n1094), .O(n1095));
  nor2   g1031(.a(n1095), .b(n962), .O(n1096));
  inv1   g1032(.a(n962), .O(n1097));
  nor2   g1033(.a(n1094), .b(n1097), .O(n1098));
  nor2   g1034(.a(n1098), .b(n1096), .O(n1099));
  inv1   g1035(.a(n1099), .O(n1100));
  nor2   g1036(.a(n1100), .b(n961), .O(n1101));
  inv1   g1037(.a(n961), .O(n1102));
  nor2   g1038(.a(n1099), .b(n1102), .O(n1103));
  nor2   g1039(.a(n1103), .b(n1101), .O(n1104));
  inv1   g1040(.a(n1104), .O(n1105));
  nor2   g1041(.a(n1105), .b(n960), .O(n1106));
  inv1   g1042(.a(n960), .O(n1107));
  nor2   g1043(.a(n1104), .b(n1107), .O(n1108));
  nor2   g1044(.a(n1108), .b(n1106), .O(n1109));
  inv1   g1045(.a(n1109), .O(G5672gat));
  inv1   g1046(.a(G511gat), .O(n1111));
  nor2   g1047(.a(n1111), .b(n65), .O(n1112));
  nor2   g1048(.a(n1106), .b(n1101), .O(n1113));
  nor2   g1049(.a(n959), .b(n68), .O(n1114));
  nor2   g1050(.a(n1096), .b(n1091), .O(n1115));
  nor2   g1051(.a(n819), .b(n82), .O(n1116));
  nor2   g1052(.a(n1086), .b(n1081), .O(n1117));
  nor2   g1053(.a(n691), .b(n104), .O(n1118));
  nor2   g1054(.a(n1076), .b(n1071), .O(n1119));
  nor2   g1055(.a(n575), .b(n138), .O(n1120));
  nor2   g1056(.a(n1066), .b(n1061), .O(n1121));
  nor2   g1057(.a(n471), .b(n184), .O(n1122));
  nor2   g1058(.a(n1056), .b(n1051), .O(n1123));
  nor2   g1059(.a(n379), .b(n242), .O(n1124));
  nor2   g1060(.a(n1046), .b(n1041), .O(n1125));
  nor2   g1061(.a(n299), .b(n312), .O(n1126));
  nor2   g1062(.a(n1036), .b(n1031), .O(n1127));
  nor2   g1063(.a(n231), .b(n394), .O(n1128));
  nor2   g1064(.a(n1026), .b(n1021), .O(n1129));
  nor2   g1065(.a(n175), .b(n488), .O(n1130));
  nor2   g1066(.a(n1016), .b(n1011), .O(n1131));
  nor2   g1067(.a(n131), .b(n594), .O(n1132));
  nor2   g1068(.a(n1006), .b(n1001), .O(n1133));
  nor2   g1069(.a(n100), .b(n712), .O(n1134));
  nor2   g1070(.a(n991), .b(n990), .O(n1135));
  nor2   g1071(.a(n1135), .b(n995), .O(n1136));
  nor2   g1072(.a(n78), .b(n842), .O(n1137));
  inv1   g1073(.a(G239gat), .O(n1138));
  nor2   g1074(.a(n66), .b(n1138), .O(n1139));
  inv1   g1075(.a(n1139), .O(n1140));
  nor2   g1076(.a(n71), .b(n984), .O(n1141));
  inv1   g1077(.a(n1141), .O(n1142));
  nor2   g1078(.a(n1142), .b(G205gat), .O(n1143));
  nor2   g1079(.a(n1143), .b(n1140), .O(n1144));
  nor2   g1080(.a(n1142), .b(n1139), .O(n1145));
  inv1   g1081(.a(n1145), .O(n1146));
  nor2   g1082(.a(n1146), .b(n843), .O(n1147));
  nor2   g1083(.a(n1147), .b(n1144), .O(n1148));
  nor2   g1084(.a(n1148), .b(n1137), .O(n1149));
  inv1   g1085(.a(n1137), .O(n1150));
  inv1   g1086(.a(n1148), .O(n1151));
  nor2   g1087(.a(n1151), .b(n1150), .O(n1152));
  nor2   g1088(.a(n1152), .b(n1149), .O(n1153));
  inv1   g1089(.a(n1153), .O(n1154));
  nor2   g1090(.a(n1154), .b(n1136), .O(n1155));
  inv1   g1091(.a(n1136), .O(n1156));
  nor2   g1092(.a(n1153), .b(n1156), .O(n1157));
  nor2   g1093(.a(n1157), .b(n1155), .O(n1158));
  inv1   g1094(.a(n1158), .O(n1159));
  nor2   g1095(.a(n1159), .b(n1134), .O(n1160));
  inv1   g1096(.a(n1134), .O(n1161));
  nor2   g1097(.a(n1158), .b(n1161), .O(n1162));
  nor2   g1098(.a(n1162), .b(n1160), .O(n1163));
  inv1   g1099(.a(n1163), .O(n1164));
  nor2   g1100(.a(n1164), .b(n1133), .O(n1165));
  inv1   g1101(.a(n1133), .O(n1166));
  nor2   g1102(.a(n1163), .b(n1166), .O(n1167));
  nor2   g1103(.a(n1167), .b(n1165), .O(n1168));
  inv1   g1104(.a(n1168), .O(n1169));
  nor2   g1105(.a(n1169), .b(n1132), .O(n1170));
  inv1   g1106(.a(n1132), .O(n1171));
  nor2   g1107(.a(n1168), .b(n1171), .O(n1172));
  nor2   g1108(.a(n1172), .b(n1170), .O(n1173));
  inv1   g1109(.a(n1173), .O(n1174));
  nor2   g1110(.a(n1174), .b(n1131), .O(n1175));
  inv1   g1111(.a(n1131), .O(n1176));
  nor2   g1112(.a(n1173), .b(n1176), .O(n1177));
  nor2   g1113(.a(n1177), .b(n1175), .O(n1178));
  inv1   g1114(.a(n1178), .O(n1179));
  nor2   g1115(.a(n1179), .b(n1130), .O(n1180));
  inv1   g1116(.a(n1130), .O(n1181));
  nor2   g1117(.a(n1178), .b(n1181), .O(n1182));
  nor2   g1118(.a(n1182), .b(n1180), .O(n1183));
  inv1   g1119(.a(n1183), .O(n1184));
  nor2   g1120(.a(n1184), .b(n1129), .O(n1185));
  inv1   g1121(.a(n1129), .O(n1186));
  nor2   g1122(.a(n1183), .b(n1186), .O(n1187));
  nor2   g1123(.a(n1187), .b(n1185), .O(n1188));
  inv1   g1124(.a(n1188), .O(n1189));
  nor2   g1125(.a(n1189), .b(n1128), .O(n1190));
  inv1   g1126(.a(n1128), .O(n1191));
  nor2   g1127(.a(n1188), .b(n1191), .O(n1192));
  nor2   g1128(.a(n1192), .b(n1190), .O(n1193));
  inv1   g1129(.a(n1193), .O(n1194));
  nor2   g1130(.a(n1194), .b(n1127), .O(n1195));
  inv1   g1131(.a(n1127), .O(n1196));
  nor2   g1132(.a(n1193), .b(n1196), .O(n1197));
  nor2   g1133(.a(n1197), .b(n1195), .O(n1198));
  inv1   g1134(.a(n1198), .O(n1199));
  nor2   g1135(.a(n1199), .b(n1126), .O(n1200));
  inv1   g1136(.a(n1126), .O(n1201));
  nor2   g1137(.a(n1198), .b(n1201), .O(n1202));
  nor2   g1138(.a(n1202), .b(n1200), .O(n1203));
  inv1   g1139(.a(n1203), .O(n1204));
  nor2   g1140(.a(n1204), .b(n1125), .O(n1205));
  inv1   g1141(.a(n1125), .O(n1206));
  nor2   g1142(.a(n1203), .b(n1206), .O(n1207));
  nor2   g1143(.a(n1207), .b(n1205), .O(n1208));
  inv1   g1144(.a(n1208), .O(n1209));
  nor2   g1145(.a(n1209), .b(n1124), .O(n1210));
  inv1   g1146(.a(n1124), .O(n1211));
  nor2   g1147(.a(n1208), .b(n1211), .O(n1212));
  nor2   g1148(.a(n1212), .b(n1210), .O(n1213));
  inv1   g1149(.a(n1213), .O(n1214));
  nor2   g1150(.a(n1214), .b(n1123), .O(n1215));
  inv1   g1151(.a(n1123), .O(n1216));
  nor2   g1152(.a(n1213), .b(n1216), .O(n1217));
  nor2   g1153(.a(n1217), .b(n1215), .O(n1218));
  inv1   g1154(.a(n1218), .O(n1219));
  nor2   g1155(.a(n1219), .b(n1122), .O(n1220));
  inv1   g1156(.a(n1122), .O(n1221));
  nor2   g1157(.a(n1218), .b(n1221), .O(n1222));
  nor2   g1158(.a(n1222), .b(n1220), .O(n1223));
  inv1   g1159(.a(n1223), .O(n1224));
  nor2   g1160(.a(n1224), .b(n1121), .O(n1225));
  inv1   g1161(.a(n1121), .O(n1226));
  nor2   g1162(.a(n1223), .b(n1226), .O(n1227));
  nor2   g1163(.a(n1227), .b(n1225), .O(n1228));
  inv1   g1164(.a(n1228), .O(n1229));
  nor2   g1165(.a(n1229), .b(n1120), .O(n1230));
  inv1   g1166(.a(n1120), .O(n1231));
  nor2   g1167(.a(n1228), .b(n1231), .O(n1232));
  nor2   g1168(.a(n1232), .b(n1230), .O(n1233));
  inv1   g1169(.a(n1233), .O(n1234));
  nor2   g1170(.a(n1234), .b(n1119), .O(n1235));
  inv1   g1171(.a(n1119), .O(n1236));
  nor2   g1172(.a(n1233), .b(n1236), .O(n1237));
  nor2   g1173(.a(n1237), .b(n1235), .O(n1238));
  inv1   g1174(.a(n1238), .O(n1239));
  nor2   g1175(.a(n1239), .b(n1118), .O(n1240));
  inv1   g1176(.a(n1118), .O(n1241));
  nor2   g1177(.a(n1238), .b(n1241), .O(n1242));
  nor2   g1178(.a(n1242), .b(n1240), .O(n1243));
  inv1   g1179(.a(n1243), .O(n1244));
  nor2   g1180(.a(n1244), .b(n1117), .O(n1245));
  inv1   g1181(.a(n1117), .O(n1246));
  nor2   g1182(.a(n1243), .b(n1246), .O(n1247));
  nor2   g1183(.a(n1247), .b(n1245), .O(n1248));
  inv1   g1184(.a(n1248), .O(n1249));
  nor2   g1185(.a(n1249), .b(n1116), .O(n1250));
  inv1   g1186(.a(n1116), .O(n1251));
  nor2   g1187(.a(n1248), .b(n1251), .O(n1252));
  nor2   g1188(.a(n1252), .b(n1250), .O(n1253));
  inv1   g1189(.a(n1253), .O(n1254));
  nor2   g1190(.a(n1254), .b(n1115), .O(n1255));
  inv1   g1191(.a(n1115), .O(n1256));
  nor2   g1192(.a(n1253), .b(n1256), .O(n1257));
  nor2   g1193(.a(n1257), .b(n1255), .O(n1258));
  inv1   g1194(.a(n1258), .O(n1259));
  nor2   g1195(.a(n1259), .b(n1114), .O(n1260));
  inv1   g1196(.a(n1114), .O(n1261));
  nor2   g1197(.a(n1258), .b(n1261), .O(n1262));
  nor2   g1198(.a(n1262), .b(n1260), .O(n1263));
  inv1   g1199(.a(n1263), .O(n1264));
  nor2   g1200(.a(n1264), .b(n1113), .O(n1265));
  inv1   g1201(.a(n1113), .O(n1266));
  nor2   g1202(.a(n1263), .b(n1266), .O(n1267));
  nor2   g1203(.a(n1267), .b(n1265), .O(n1268));
  inv1   g1204(.a(n1268), .O(n1269));
  nor2   g1205(.a(n1269), .b(n1112), .O(n1270));
  inv1   g1206(.a(n1112), .O(n1271));
  nor2   g1207(.a(n1268), .b(n1271), .O(n1272));
  nor2   g1208(.a(n1272), .b(n1270), .O(n1273));
  inv1   g1209(.a(n1273), .O(G5971gat));
  inv1   g1210(.a(G528gat), .O(n1275));
  nor2   g1211(.a(n1275), .b(n65), .O(n1276));
  nor2   g1212(.a(n1270), .b(n1265), .O(n1277));
  nor2   g1213(.a(n1111), .b(n68), .O(n1278));
  nor2   g1214(.a(n1260), .b(n1255), .O(n1279));
  nor2   g1215(.a(n959), .b(n82), .O(n1280));
  nor2   g1216(.a(n1250), .b(n1245), .O(n1281));
  nor2   g1217(.a(n819), .b(n104), .O(n1282));
  nor2   g1218(.a(n1240), .b(n1235), .O(n1283));
  nor2   g1219(.a(n691), .b(n138), .O(n1284));
  nor2   g1220(.a(n1230), .b(n1225), .O(n1285));
  nor2   g1221(.a(n575), .b(n184), .O(n1286));
  nor2   g1222(.a(n1220), .b(n1215), .O(n1287));
  nor2   g1223(.a(n471), .b(n242), .O(n1288));
  nor2   g1224(.a(n1210), .b(n1205), .O(n1289));
  nor2   g1225(.a(n379), .b(n312), .O(n1290));
  nor2   g1226(.a(n1200), .b(n1195), .O(n1291));
  nor2   g1227(.a(n299), .b(n394), .O(n1292));
  nor2   g1228(.a(n1190), .b(n1185), .O(n1293));
  nor2   g1229(.a(n231), .b(n488), .O(n1294));
  nor2   g1230(.a(n1180), .b(n1175), .O(n1295));
  nor2   g1231(.a(n175), .b(n594), .O(n1296));
  nor2   g1232(.a(n1170), .b(n1165), .O(n1297));
  nor2   g1233(.a(n131), .b(n712), .O(n1298));
  nor2   g1234(.a(n1160), .b(n1155), .O(n1299));
  nor2   g1235(.a(n100), .b(n842), .O(n1300));
  nor2   g1236(.a(n1145), .b(n1144), .O(n1301));
  nor2   g1237(.a(n1301), .b(n1149), .O(n1302));
  nor2   g1238(.a(n78), .b(n984), .O(n1303));
  inv1   g1239(.a(G256gat), .O(n1304));
  nor2   g1240(.a(n66), .b(n1304), .O(n1305));
  inv1   g1241(.a(n1305), .O(n1306));
  nor2   g1242(.a(n71), .b(n1138), .O(n1307));
  inv1   g1243(.a(n1307), .O(n1308));
  nor2   g1244(.a(n1308), .b(G222gat), .O(n1309));
  nor2   g1245(.a(n1309), .b(n1306), .O(n1310));
  nor2   g1246(.a(n1308), .b(n1305), .O(n1311));
  inv1   g1247(.a(n1311), .O(n1312));
  nor2   g1248(.a(n1312), .b(n985), .O(n1313));
  nor2   g1249(.a(n1313), .b(n1310), .O(n1314));
  nor2   g1250(.a(n1314), .b(n1303), .O(n1315));
  inv1   g1251(.a(n1303), .O(n1316));
  inv1   g1252(.a(n1314), .O(n1317));
  nor2   g1253(.a(n1317), .b(n1316), .O(n1318));
  nor2   g1254(.a(n1318), .b(n1315), .O(n1319));
  inv1   g1255(.a(n1319), .O(n1320));
  nor2   g1256(.a(n1320), .b(n1302), .O(n1321));
  inv1   g1257(.a(n1302), .O(n1322));
  nor2   g1258(.a(n1319), .b(n1322), .O(n1323));
  nor2   g1259(.a(n1323), .b(n1321), .O(n1324));
  inv1   g1260(.a(n1324), .O(n1325));
  nor2   g1261(.a(n1325), .b(n1300), .O(n1326));
  inv1   g1262(.a(n1300), .O(n1327));
  nor2   g1263(.a(n1324), .b(n1327), .O(n1328));
  nor2   g1264(.a(n1328), .b(n1326), .O(n1329));
  inv1   g1265(.a(n1329), .O(n1330));
  nor2   g1266(.a(n1330), .b(n1299), .O(n1331));
  inv1   g1267(.a(n1299), .O(n1332));
  nor2   g1268(.a(n1329), .b(n1332), .O(n1333));
  nor2   g1269(.a(n1333), .b(n1331), .O(n1334));
  inv1   g1270(.a(n1334), .O(n1335));
  nor2   g1271(.a(n1335), .b(n1298), .O(n1336));
  inv1   g1272(.a(n1298), .O(n1337));
  nor2   g1273(.a(n1334), .b(n1337), .O(n1338));
  nor2   g1274(.a(n1338), .b(n1336), .O(n1339));
  inv1   g1275(.a(n1339), .O(n1340));
  nor2   g1276(.a(n1340), .b(n1297), .O(n1341));
  inv1   g1277(.a(n1297), .O(n1342));
  nor2   g1278(.a(n1339), .b(n1342), .O(n1343));
  nor2   g1279(.a(n1343), .b(n1341), .O(n1344));
  inv1   g1280(.a(n1344), .O(n1345));
  nor2   g1281(.a(n1345), .b(n1296), .O(n1346));
  inv1   g1282(.a(n1296), .O(n1347));
  nor2   g1283(.a(n1344), .b(n1347), .O(n1348));
  nor2   g1284(.a(n1348), .b(n1346), .O(n1349));
  inv1   g1285(.a(n1349), .O(n1350));
  nor2   g1286(.a(n1350), .b(n1295), .O(n1351));
  inv1   g1287(.a(n1295), .O(n1352));
  nor2   g1288(.a(n1349), .b(n1352), .O(n1353));
  nor2   g1289(.a(n1353), .b(n1351), .O(n1354));
  inv1   g1290(.a(n1354), .O(n1355));
  nor2   g1291(.a(n1355), .b(n1294), .O(n1356));
  inv1   g1292(.a(n1294), .O(n1357));
  nor2   g1293(.a(n1354), .b(n1357), .O(n1358));
  nor2   g1294(.a(n1358), .b(n1356), .O(n1359));
  inv1   g1295(.a(n1359), .O(n1360));
  nor2   g1296(.a(n1360), .b(n1293), .O(n1361));
  inv1   g1297(.a(n1293), .O(n1362));
  nor2   g1298(.a(n1359), .b(n1362), .O(n1363));
  nor2   g1299(.a(n1363), .b(n1361), .O(n1364));
  inv1   g1300(.a(n1364), .O(n1365));
  nor2   g1301(.a(n1365), .b(n1292), .O(n1366));
  inv1   g1302(.a(n1292), .O(n1367));
  nor2   g1303(.a(n1364), .b(n1367), .O(n1368));
  nor2   g1304(.a(n1368), .b(n1366), .O(n1369));
  inv1   g1305(.a(n1369), .O(n1370));
  nor2   g1306(.a(n1370), .b(n1291), .O(n1371));
  inv1   g1307(.a(n1291), .O(n1372));
  nor2   g1308(.a(n1369), .b(n1372), .O(n1373));
  nor2   g1309(.a(n1373), .b(n1371), .O(n1374));
  inv1   g1310(.a(n1374), .O(n1375));
  nor2   g1311(.a(n1375), .b(n1290), .O(n1376));
  inv1   g1312(.a(n1290), .O(n1377));
  nor2   g1313(.a(n1374), .b(n1377), .O(n1378));
  nor2   g1314(.a(n1378), .b(n1376), .O(n1379));
  inv1   g1315(.a(n1379), .O(n1380));
  nor2   g1316(.a(n1380), .b(n1289), .O(n1381));
  inv1   g1317(.a(n1289), .O(n1382));
  nor2   g1318(.a(n1379), .b(n1382), .O(n1383));
  nor2   g1319(.a(n1383), .b(n1381), .O(n1384));
  inv1   g1320(.a(n1384), .O(n1385));
  nor2   g1321(.a(n1385), .b(n1288), .O(n1386));
  inv1   g1322(.a(n1288), .O(n1387));
  nor2   g1323(.a(n1384), .b(n1387), .O(n1388));
  nor2   g1324(.a(n1388), .b(n1386), .O(n1389));
  inv1   g1325(.a(n1389), .O(n1390));
  nor2   g1326(.a(n1390), .b(n1287), .O(n1391));
  inv1   g1327(.a(n1287), .O(n1392));
  nor2   g1328(.a(n1389), .b(n1392), .O(n1393));
  nor2   g1329(.a(n1393), .b(n1391), .O(n1394));
  inv1   g1330(.a(n1394), .O(n1395));
  nor2   g1331(.a(n1395), .b(n1286), .O(n1396));
  inv1   g1332(.a(n1286), .O(n1397));
  nor2   g1333(.a(n1394), .b(n1397), .O(n1398));
  nor2   g1334(.a(n1398), .b(n1396), .O(n1399));
  inv1   g1335(.a(n1399), .O(n1400));
  nor2   g1336(.a(n1400), .b(n1285), .O(n1401));
  inv1   g1337(.a(n1285), .O(n1402));
  nor2   g1338(.a(n1399), .b(n1402), .O(n1403));
  nor2   g1339(.a(n1403), .b(n1401), .O(n1404));
  inv1   g1340(.a(n1404), .O(n1405));
  nor2   g1341(.a(n1405), .b(n1284), .O(n1406));
  inv1   g1342(.a(n1284), .O(n1407));
  nor2   g1343(.a(n1404), .b(n1407), .O(n1408));
  nor2   g1344(.a(n1408), .b(n1406), .O(n1409));
  inv1   g1345(.a(n1409), .O(n1410));
  nor2   g1346(.a(n1410), .b(n1283), .O(n1411));
  inv1   g1347(.a(n1283), .O(n1412));
  nor2   g1348(.a(n1409), .b(n1412), .O(n1413));
  nor2   g1349(.a(n1413), .b(n1411), .O(n1414));
  inv1   g1350(.a(n1414), .O(n1415));
  nor2   g1351(.a(n1415), .b(n1282), .O(n1416));
  inv1   g1352(.a(n1282), .O(n1417));
  nor2   g1353(.a(n1414), .b(n1417), .O(n1418));
  nor2   g1354(.a(n1418), .b(n1416), .O(n1419));
  inv1   g1355(.a(n1419), .O(n1420));
  nor2   g1356(.a(n1420), .b(n1281), .O(n1421));
  inv1   g1357(.a(n1281), .O(n1422));
  nor2   g1358(.a(n1419), .b(n1422), .O(n1423));
  nor2   g1359(.a(n1423), .b(n1421), .O(n1424));
  inv1   g1360(.a(n1424), .O(n1425));
  nor2   g1361(.a(n1425), .b(n1280), .O(n1426));
  inv1   g1362(.a(n1280), .O(n1427));
  nor2   g1363(.a(n1424), .b(n1427), .O(n1428));
  nor2   g1364(.a(n1428), .b(n1426), .O(n1429));
  inv1   g1365(.a(n1429), .O(n1430));
  nor2   g1366(.a(n1430), .b(n1279), .O(n1431));
  inv1   g1367(.a(n1279), .O(n1432));
  nor2   g1368(.a(n1429), .b(n1432), .O(n1433));
  nor2   g1369(.a(n1433), .b(n1431), .O(n1434));
  inv1   g1370(.a(n1434), .O(n1435));
  nor2   g1371(.a(n1435), .b(n1278), .O(n1436));
  inv1   g1372(.a(n1278), .O(n1437));
  nor2   g1373(.a(n1434), .b(n1437), .O(n1438));
  nor2   g1374(.a(n1438), .b(n1436), .O(n1439));
  inv1   g1375(.a(n1439), .O(n1440));
  nor2   g1376(.a(n1440), .b(n1277), .O(n1441));
  inv1   g1377(.a(n1277), .O(n1442));
  nor2   g1378(.a(n1439), .b(n1442), .O(n1443));
  nor2   g1379(.a(n1443), .b(n1441), .O(n1444));
  inv1   g1380(.a(n1444), .O(n1445));
  nor2   g1381(.a(n1445), .b(n1276), .O(n1446));
  inv1   g1382(.a(n1276), .O(n1447));
  nor2   g1383(.a(n1444), .b(n1447), .O(n1448));
  nor2   g1384(.a(n1448), .b(n1446), .O(n1449));
  inv1   g1385(.a(n1449), .O(G6123gat));
  nor2   g1386(.a(n1446), .b(n1441), .O(n1451));
  nor2   g1387(.a(n1275), .b(n68), .O(n1452));
  nor2   g1388(.a(n1436), .b(n1431), .O(n1453));
  nor2   g1389(.a(n1111), .b(n82), .O(n1454));
  nor2   g1390(.a(n1426), .b(n1421), .O(n1455));
  nor2   g1391(.a(n959), .b(n104), .O(n1456));
  nor2   g1392(.a(n1416), .b(n1411), .O(n1457));
  nor2   g1393(.a(n819), .b(n138), .O(n1458));
  nor2   g1394(.a(n1406), .b(n1401), .O(n1459));
  nor2   g1395(.a(n691), .b(n184), .O(n1460));
  nor2   g1396(.a(n1396), .b(n1391), .O(n1461));
  nor2   g1397(.a(n575), .b(n242), .O(n1462));
  nor2   g1398(.a(n1386), .b(n1381), .O(n1463));
  nor2   g1399(.a(n471), .b(n312), .O(n1464));
  nor2   g1400(.a(n1376), .b(n1371), .O(n1465));
  nor2   g1401(.a(n379), .b(n394), .O(n1466));
  nor2   g1402(.a(n1366), .b(n1361), .O(n1467));
  nor2   g1403(.a(n299), .b(n488), .O(n1468));
  nor2   g1404(.a(n1356), .b(n1351), .O(n1469));
  nor2   g1405(.a(n231), .b(n594), .O(n1470));
  nor2   g1406(.a(n1346), .b(n1341), .O(n1471));
  nor2   g1407(.a(n175), .b(n712), .O(n1472));
  nor2   g1408(.a(n1336), .b(n1331), .O(n1473));
  nor2   g1409(.a(n131), .b(n842), .O(n1474));
  nor2   g1410(.a(n1326), .b(n1321), .O(n1475));
  nor2   g1411(.a(n100), .b(n984), .O(n1476));
  nor2   g1412(.a(n1311), .b(n1310), .O(n1477));
  nor2   g1413(.a(n1477), .b(n1315), .O(n1478));
  nor2   g1414(.a(n78), .b(n1138), .O(n1479));
  nor2   g1415(.a(n71), .b(n1304), .O(n1480));
  inv1   g1416(.a(n1480), .O(n1481));
  nor2   g1417(.a(n1481), .b(n1139), .O(n1482));
  inv1   g1418(.a(n1482), .O(n1483));
  nor2   g1419(.a(n1483), .b(n1479), .O(n1484));
  inv1   g1420(.a(n1479), .O(n1485));
  nor2   g1421(.a(n1482), .b(n1485), .O(n1486));
  nor2   g1422(.a(n1486), .b(n1484), .O(n1487));
  inv1   g1423(.a(n1487), .O(n1488));
  nor2   g1424(.a(n1488), .b(n1478), .O(n1489));
  inv1   g1425(.a(n1478), .O(n1490));
  nor2   g1426(.a(n1487), .b(n1490), .O(n1491));
  nor2   g1427(.a(n1491), .b(n1489), .O(n1492));
  inv1   g1428(.a(n1492), .O(n1493));
  nor2   g1429(.a(n1493), .b(n1476), .O(n1494));
  inv1   g1430(.a(n1476), .O(n1495));
  nor2   g1431(.a(n1492), .b(n1495), .O(n1496));
  nor2   g1432(.a(n1496), .b(n1494), .O(n1497));
  inv1   g1433(.a(n1497), .O(n1498));
  nor2   g1434(.a(n1498), .b(n1475), .O(n1499));
  inv1   g1435(.a(n1475), .O(n1500));
  nor2   g1436(.a(n1497), .b(n1500), .O(n1501));
  nor2   g1437(.a(n1501), .b(n1499), .O(n1502));
  inv1   g1438(.a(n1502), .O(n1503));
  nor2   g1439(.a(n1503), .b(n1474), .O(n1504));
  inv1   g1440(.a(n1474), .O(n1505));
  nor2   g1441(.a(n1502), .b(n1505), .O(n1506));
  nor2   g1442(.a(n1506), .b(n1504), .O(n1507));
  inv1   g1443(.a(n1507), .O(n1508));
  nor2   g1444(.a(n1508), .b(n1473), .O(n1509));
  inv1   g1445(.a(n1473), .O(n1510));
  nor2   g1446(.a(n1507), .b(n1510), .O(n1511));
  nor2   g1447(.a(n1511), .b(n1509), .O(n1512));
  inv1   g1448(.a(n1512), .O(n1513));
  nor2   g1449(.a(n1513), .b(n1472), .O(n1514));
  inv1   g1450(.a(n1472), .O(n1515));
  nor2   g1451(.a(n1512), .b(n1515), .O(n1516));
  nor2   g1452(.a(n1516), .b(n1514), .O(n1517));
  inv1   g1453(.a(n1517), .O(n1518));
  nor2   g1454(.a(n1518), .b(n1471), .O(n1519));
  inv1   g1455(.a(n1471), .O(n1520));
  nor2   g1456(.a(n1517), .b(n1520), .O(n1521));
  nor2   g1457(.a(n1521), .b(n1519), .O(n1522));
  inv1   g1458(.a(n1522), .O(n1523));
  nor2   g1459(.a(n1523), .b(n1470), .O(n1524));
  inv1   g1460(.a(n1470), .O(n1525));
  nor2   g1461(.a(n1522), .b(n1525), .O(n1526));
  nor2   g1462(.a(n1526), .b(n1524), .O(n1527));
  inv1   g1463(.a(n1527), .O(n1528));
  nor2   g1464(.a(n1528), .b(n1469), .O(n1529));
  inv1   g1465(.a(n1469), .O(n1530));
  nor2   g1466(.a(n1527), .b(n1530), .O(n1531));
  nor2   g1467(.a(n1531), .b(n1529), .O(n1532));
  inv1   g1468(.a(n1532), .O(n1533));
  nor2   g1469(.a(n1533), .b(n1468), .O(n1534));
  inv1   g1470(.a(n1468), .O(n1535));
  nor2   g1471(.a(n1532), .b(n1535), .O(n1536));
  nor2   g1472(.a(n1536), .b(n1534), .O(n1537));
  inv1   g1473(.a(n1537), .O(n1538));
  nor2   g1474(.a(n1538), .b(n1467), .O(n1539));
  inv1   g1475(.a(n1467), .O(n1540));
  nor2   g1476(.a(n1537), .b(n1540), .O(n1541));
  nor2   g1477(.a(n1541), .b(n1539), .O(n1542));
  inv1   g1478(.a(n1542), .O(n1543));
  nor2   g1479(.a(n1543), .b(n1466), .O(n1544));
  inv1   g1480(.a(n1466), .O(n1545));
  nor2   g1481(.a(n1542), .b(n1545), .O(n1546));
  nor2   g1482(.a(n1546), .b(n1544), .O(n1547));
  inv1   g1483(.a(n1547), .O(n1548));
  nor2   g1484(.a(n1548), .b(n1465), .O(n1549));
  inv1   g1485(.a(n1465), .O(n1550));
  nor2   g1486(.a(n1547), .b(n1550), .O(n1551));
  nor2   g1487(.a(n1551), .b(n1549), .O(n1552));
  inv1   g1488(.a(n1552), .O(n1553));
  nor2   g1489(.a(n1553), .b(n1464), .O(n1554));
  inv1   g1490(.a(n1464), .O(n1555));
  nor2   g1491(.a(n1552), .b(n1555), .O(n1556));
  nor2   g1492(.a(n1556), .b(n1554), .O(n1557));
  inv1   g1493(.a(n1557), .O(n1558));
  nor2   g1494(.a(n1558), .b(n1463), .O(n1559));
  inv1   g1495(.a(n1463), .O(n1560));
  nor2   g1496(.a(n1557), .b(n1560), .O(n1561));
  nor2   g1497(.a(n1561), .b(n1559), .O(n1562));
  inv1   g1498(.a(n1562), .O(n1563));
  nor2   g1499(.a(n1563), .b(n1462), .O(n1564));
  inv1   g1500(.a(n1462), .O(n1565));
  nor2   g1501(.a(n1562), .b(n1565), .O(n1566));
  nor2   g1502(.a(n1566), .b(n1564), .O(n1567));
  inv1   g1503(.a(n1567), .O(n1568));
  nor2   g1504(.a(n1568), .b(n1461), .O(n1569));
  inv1   g1505(.a(n1461), .O(n1570));
  nor2   g1506(.a(n1567), .b(n1570), .O(n1571));
  nor2   g1507(.a(n1571), .b(n1569), .O(n1572));
  inv1   g1508(.a(n1572), .O(n1573));
  nor2   g1509(.a(n1573), .b(n1460), .O(n1574));
  inv1   g1510(.a(n1460), .O(n1575));
  nor2   g1511(.a(n1572), .b(n1575), .O(n1576));
  nor2   g1512(.a(n1576), .b(n1574), .O(n1577));
  inv1   g1513(.a(n1577), .O(n1578));
  nor2   g1514(.a(n1578), .b(n1459), .O(n1579));
  inv1   g1515(.a(n1459), .O(n1580));
  nor2   g1516(.a(n1577), .b(n1580), .O(n1581));
  nor2   g1517(.a(n1581), .b(n1579), .O(n1582));
  inv1   g1518(.a(n1582), .O(n1583));
  nor2   g1519(.a(n1583), .b(n1458), .O(n1584));
  inv1   g1520(.a(n1458), .O(n1585));
  nor2   g1521(.a(n1582), .b(n1585), .O(n1586));
  nor2   g1522(.a(n1586), .b(n1584), .O(n1587));
  inv1   g1523(.a(n1587), .O(n1588));
  nor2   g1524(.a(n1588), .b(n1457), .O(n1589));
  inv1   g1525(.a(n1457), .O(n1590));
  nor2   g1526(.a(n1587), .b(n1590), .O(n1591));
  nor2   g1527(.a(n1591), .b(n1589), .O(n1592));
  inv1   g1528(.a(n1592), .O(n1593));
  nor2   g1529(.a(n1593), .b(n1456), .O(n1594));
  inv1   g1530(.a(n1456), .O(n1595));
  nor2   g1531(.a(n1592), .b(n1595), .O(n1596));
  nor2   g1532(.a(n1596), .b(n1594), .O(n1597));
  inv1   g1533(.a(n1597), .O(n1598));
  nor2   g1534(.a(n1598), .b(n1455), .O(n1599));
  inv1   g1535(.a(n1455), .O(n1600));
  nor2   g1536(.a(n1597), .b(n1600), .O(n1601));
  nor2   g1537(.a(n1601), .b(n1599), .O(n1602));
  inv1   g1538(.a(n1602), .O(n1603));
  nor2   g1539(.a(n1603), .b(n1454), .O(n1604));
  inv1   g1540(.a(n1454), .O(n1605));
  nor2   g1541(.a(n1602), .b(n1605), .O(n1606));
  nor2   g1542(.a(n1606), .b(n1604), .O(n1607));
  inv1   g1543(.a(n1607), .O(n1608));
  nor2   g1544(.a(n1608), .b(n1453), .O(n1609));
  inv1   g1545(.a(n1453), .O(n1610));
  nor2   g1546(.a(n1607), .b(n1610), .O(n1611));
  nor2   g1547(.a(n1611), .b(n1609), .O(n1612));
  inv1   g1548(.a(n1612), .O(n1613));
  nor2   g1549(.a(n1613), .b(n1452), .O(n1614));
  inv1   g1550(.a(n1452), .O(n1615));
  nor2   g1551(.a(n1612), .b(n1615), .O(n1616));
  nor2   g1552(.a(n1616), .b(n1614), .O(n1617));
  inv1   g1553(.a(n1617), .O(n1618));
  nor2   g1554(.a(n1618), .b(n1451), .O(n1619));
  inv1   g1555(.a(n1451), .O(n1620));
  nor2   g1556(.a(n1617), .b(n1620), .O(n1621));
  nor2   g1557(.a(n1621), .b(n1619), .O(G6150gat));
  nor2   g1558(.a(n1614), .b(n1609), .O(n1623));
  nor2   g1559(.a(n1275), .b(n82), .O(n1624));
  nor2   g1560(.a(n1604), .b(n1599), .O(n1625));
  nor2   g1561(.a(n1111), .b(n104), .O(n1626));
  nor2   g1562(.a(n1594), .b(n1589), .O(n1627));
  nor2   g1563(.a(n959), .b(n138), .O(n1628));
  nor2   g1564(.a(n1584), .b(n1579), .O(n1629));
  nor2   g1565(.a(n819), .b(n184), .O(n1630));
  nor2   g1566(.a(n1574), .b(n1569), .O(n1631));
  nor2   g1567(.a(n691), .b(n242), .O(n1632));
  nor2   g1568(.a(n1564), .b(n1559), .O(n1633));
  nor2   g1569(.a(n575), .b(n312), .O(n1634));
  nor2   g1570(.a(n1554), .b(n1549), .O(n1635));
  nor2   g1571(.a(n471), .b(n394), .O(n1636));
  nor2   g1572(.a(n1544), .b(n1539), .O(n1637));
  nor2   g1573(.a(n379), .b(n488), .O(n1638));
  nor2   g1574(.a(n1534), .b(n1529), .O(n1639));
  nor2   g1575(.a(n299), .b(n594), .O(n1640));
  nor2   g1576(.a(n1524), .b(n1519), .O(n1641));
  nor2   g1577(.a(n231), .b(n712), .O(n1642));
  nor2   g1578(.a(n1514), .b(n1509), .O(n1643));
  nor2   g1579(.a(n175), .b(n842), .O(n1644));
  nor2   g1580(.a(n1504), .b(n1499), .O(n1645));
  nor2   g1581(.a(n131), .b(n984), .O(n1646));
  nor2   g1582(.a(n1494), .b(n1489), .O(n1647));
  nor2   g1583(.a(n100), .b(n1138), .O(n1648));
  nor2   g1584(.a(n1308), .b(n66), .O(n1649));
  nor2   g1585(.a(n1649), .b(G307gat), .O(n1650));
  nor2   g1586(.a(n1650), .b(n1304), .O(n1651));
  inv1   g1587(.a(n1651), .O(n1652));
  nor2   g1588(.a(n1485), .b(n71), .O(n1653));
  nor2   g1589(.a(n1653), .b(n1652), .O(n1654));
  inv1   g1590(.a(n1654), .O(n1655));
  nor2   g1591(.a(n1655), .b(n1648), .O(n1656));
  inv1   g1592(.a(n1648), .O(n1657));
  nor2   g1593(.a(n1654), .b(n1657), .O(n1658));
  nor2   g1594(.a(n1658), .b(n1656), .O(n1659));
  inv1   g1595(.a(n1659), .O(n1660));
  nor2   g1596(.a(n1660), .b(n1647), .O(n1661));
  inv1   g1597(.a(n1647), .O(n1662));
  nor2   g1598(.a(n1659), .b(n1662), .O(n1663));
  nor2   g1599(.a(n1663), .b(n1661), .O(n1664));
  inv1   g1600(.a(n1664), .O(n1665));
  nor2   g1601(.a(n1665), .b(n1646), .O(n1666));
  inv1   g1602(.a(n1646), .O(n1667));
  nor2   g1603(.a(n1664), .b(n1667), .O(n1668));
  nor2   g1604(.a(n1668), .b(n1666), .O(n1669));
  inv1   g1605(.a(n1669), .O(n1670));
  nor2   g1606(.a(n1670), .b(n1645), .O(n1671));
  inv1   g1607(.a(n1645), .O(n1672));
  nor2   g1608(.a(n1669), .b(n1672), .O(n1673));
  nor2   g1609(.a(n1673), .b(n1671), .O(n1674));
  inv1   g1610(.a(n1674), .O(n1675));
  nor2   g1611(.a(n1675), .b(n1644), .O(n1676));
  inv1   g1612(.a(n1644), .O(n1677));
  nor2   g1613(.a(n1674), .b(n1677), .O(n1678));
  nor2   g1614(.a(n1678), .b(n1676), .O(n1679));
  inv1   g1615(.a(n1679), .O(n1680));
  nor2   g1616(.a(n1680), .b(n1643), .O(n1681));
  inv1   g1617(.a(n1643), .O(n1682));
  nor2   g1618(.a(n1679), .b(n1682), .O(n1683));
  nor2   g1619(.a(n1683), .b(n1681), .O(n1684));
  inv1   g1620(.a(n1684), .O(n1685));
  nor2   g1621(.a(n1685), .b(n1642), .O(n1686));
  inv1   g1622(.a(n1642), .O(n1687));
  nor2   g1623(.a(n1684), .b(n1687), .O(n1688));
  nor2   g1624(.a(n1688), .b(n1686), .O(n1689));
  inv1   g1625(.a(n1689), .O(n1690));
  nor2   g1626(.a(n1690), .b(n1641), .O(n1691));
  inv1   g1627(.a(n1641), .O(n1692));
  nor2   g1628(.a(n1689), .b(n1692), .O(n1693));
  nor2   g1629(.a(n1693), .b(n1691), .O(n1694));
  inv1   g1630(.a(n1694), .O(n1695));
  nor2   g1631(.a(n1695), .b(n1640), .O(n1696));
  inv1   g1632(.a(n1640), .O(n1697));
  nor2   g1633(.a(n1694), .b(n1697), .O(n1698));
  nor2   g1634(.a(n1698), .b(n1696), .O(n1699));
  inv1   g1635(.a(n1699), .O(n1700));
  nor2   g1636(.a(n1700), .b(n1639), .O(n1701));
  inv1   g1637(.a(n1639), .O(n1702));
  nor2   g1638(.a(n1699), .b(n1702), .O(n1703));
  nor2   g1639(.a(n1703), .b(n1701), .O(n1704));
  inv1   g1640(.a(n1704), .O(n1705));
  nor2   g1641(.a(n1705), .b(n1638), .O(n1706));
  inv1   g1642(.a(n1638), .O(n1707));
  nor2   g1643(.a(n1704), .b(n1707), .O(n1708));
  nor2   g1644(.a(n1708), .b(n1706), .O(n1709));
  inv1   g1645(.a(n1709), .O(n1710));
  nor2   g1646(.a(n1710), .b(n1637), .O(n1711));
  inv1   g1647(.a(n1637), .O(n1712));
  nor2   g1648(.a(n1709), .b(n1712), .O(n1713));
  nor2   g1649(.a(n1713), .b(n1711), .O(n1714));
  inv1   g1650(.a(n1714), .O(n1715));
  nor2   g1651(.a(n1715), .b(n1636), .O(n1716));
  inv1   g1652(.a(n1636), .O(n1717));
  nor2   g1653(.a(n1714), .b(n1717), .O(n1718));
  nor2   g1654(.a(n1718), .b(n1716), .O(n1719));
  inv1   g1655(.a(n1719), .O(n1720));
  nor2   g1656(.a(n1720), .b(n1635), .O(n1721));
  inv1   g1657(.a(n1635), .O(n1722));
  nor2   g1658(.a(n1719), .b(n1722), .O(n1723));
  nor2   g1659(.a(n1723), .b(n1721), .O(n1724));
  inv1   g1660(.a(n1724), .O(n1725));
  nor2   g1661(.a(n1725), .b(n1634), .O(n1726));
  inv1   g1662(.a(n1634), .O(n1727));
  nor2   g1663(.a(n1724), .b(n1727), .O(n1728));
  nor2   g1664(.a(n1728), .b(n1726), .O(n1729));
  inv1   g1665(.a(n1729), .O(n1730));
  nor2   g1666(.a(n1730), .b(n1633), .O(n1731));
  inv1   g1667(.a(n1633), .O(n1732));
  nor2   g1668(.a(n1729), .b(n1732), .O(n1733));
  nor2   g1669(.a(n1733), .b(n1731), .O(n1734));
  inv1   g1670(.a(n1734), .O(n1735));
  nor2   g1671(.a(n1735), .b(n1632), .O(n1736));
  inv1   g1672(.a(n1632), .O(n1737));
  nor2   g1673(.a(n1734), .b(n1737), .O(n1738));
  nor2   g1674(.a(n1738), .b(n1736), .O(n1739));
  inv1   g1675(.a(n1739), .O(n1740));
  nor2   g1676(.a(n1740), .b(n1631), .O(n1741));
  inv1   g1677(.a(n1631), .O(n1742));
  nor2   g1678(.a(n1739), .b(n1742), .O(n1743));
  nor2   g1679(.a(n1743), .b(n1741), .O(n1744));
  inv1   g1680(.a(n1744), .O(n1745));
  nor2   g1681(.a(n1745), .b(n1630), .O(n1746));
  inv1   g1682(.a(n1630), .O(n1747));
  nor2   g1683(.a(n1744), .b(n1747), .O(n1748));
  nor2   g1684(.a(n1748), .b(n1746), .O(n1749));
  inv1   g1685(.a(n1749), .O(n1750));
  nor2   g1686(.a(n1750), .b(n1629), .O(n1751));
  inv1   g1687(.a(n1629), .O(n1752));
  nor2   g1688(.a(n1749), .b(n1752), .O(n1753));
  nor2   g1689(.a(n1753), .b(n1751), .O(n1754));
  inv1   g1690(.a(n1754), .O(n1755));
  nor2   g1691(.a(n1755), .b(n1628), .O(n1756));
  inv1   g1692(.a(n1628), .O(n1757));
  nor2   g1693(.a(n1754), .b(n1757), .O(n1758));
  nor2   g1694(.a(n1758), .b(n1756), .O(n1759));
  inv1   g1695(.a(n1759), .O(n1760));
  nor2   g1696(.a(n1760), .b(n1627), .O(n1761));
  inv1   g1697(.a(n1627), .O(n1762));
  nor2   g1698(.a(n1759), .b(n1762), .O(n1763));
  nor2   g1699(.a(n1763), .b(n1761), .O(n1764));
  inv1   g1700(.a(n1764), .O(n1765));
  nor2   g1701(.a(n1765), .b(n1626), .O(n1766));
  inv1   g1702(.a(n1626), .O(n1767));
  nor2   g1703(.a(n1764), .b(n1767), .O(n1768));
  nor2   g1704(.a(n1768), .b(n1766), .O(n1769));
  inv1   g1705(.a(n1769), .O(n1770));
  nor2   g1706(.a(n1770), .b(n1625), .O(n1771));
  inv1   g1707(.a(n1625), .O(n1772));
  nor2   g1708(.a(n1769), .b(n1772), .O(n1773));
  nor2   g1709(.a(n1773), .b(n1771), .O(n1774));
  inv1   g1710(.a(n1774), .O(n1775));
  nor2   g1711(.a(n1775), .b(n1624), .O(n1776));
  inv1   g1712(.a(n1624), .O(n1777));
  nor2   g1713(.a(n1774), .b(n1777), .O(n1778));
  nor2   g1714(.a(n1778), .b(n1776), .O(n1779));
  inv1   g1715(.a(n1779), .O(n1780));
  nor2   g1716(.a(n1780), .b(n1623), .O(n1781));
  inv1   g1717(.a(n1623), .O(n1782));
  nor2   g1718(.a(n1779), .b(n1782), .O(n1783));
  nor2   g1719(.a(n1783), .b(n1781), .O(n1784));
  inv1   g1720(.a(n1784), .O(n1785));
  nor2   g1721(.a(n1785), .b(n1621), .O(n1786));
  inv1   g1722(.a(n1621), .O(n1787));
  nor2   g1723(.a(n1784), .b(n1787), .O(n1788));
  nor2   g1724(.a(n1788), .b(n1786), .O(n1789));
  inv1   g1725(.a(n1789), .O(G6160gat));
  nor2   g1726(.a(n1786), .b(n1781), .O(n1791));
  nor2   g1727(.a(n1776), .b(n1771), .O(n1792));
  nor2   g1728(.a(n1275), .b(n104), .O(n1793));
  nor2   g1729(.a(n1766), .b(n1761), .O(n1794));
  nor2   g1730(.a(n1111), .b(n138), .O(n1795));
  nor2   g1731(.a(n1756), .b(n1751), .O(n1796));
  nor2   g1732(.a(n959), .b(n184), .O(n1797));
  nor2   g1733(.a(n1746), .b(n1741), .O(n1798));
  nor2   g1734(.a(n819), .b(n242), .O(n1799));
  nor2   g1735(.a(n1736), .b(n1731), .O(n1800));
  nor2   g1736(.a(n691), .b(n312), .O(n1801));
  nor2   g1737(.a(n1726), .b(n1721), .O(n1802));
  nor2   g1738(.a(n575), .b(n394), .O(n1803));
  nor2   g1739(.a(n1716), .b(n1711), .O(n1804));
  nor2   g1740(.a(n471), .b(n488), .O(n1805));
  nor2   g1741(.a(n1706), .b(n1701), .O(n1806));
  nor2   g1742(.a(n379), .b(n594), .O(n1807));
  nor2   g1743(.a(n1696), .b(n1691), .O(n1808));
  nor2   g1744(.a(n299), .b(n712), .O(n1809));
  nor2   g1745(.a(n1686), .b(n1681), .O(n1810));
  nor2   g1746(.a(n231), .b(n842), .O(n1811));
  nor2   g1747(.a(n1676), .b(n1671), .O(n1812));
  nor2   g1748(.a(n175), .b(n984), .O(n1813));
  nor2   g1749(.a(n1666), .b(n1661), .O(n1814));
  nor2   g1750(.a(n131), .b(n1138), .O(n1815));
  nor2   g1751(.a(n100), .b(n1304), .O(n1816));
  nor2   g1752(.a(n1656), .b(n1652), .O(n1817));
  nor2   g1753(.a(n1817), .b(n1816), .O(n1818));
  inv1   g1754(.a(n1817), .O(n1819));
  nor2   g1755(.a(n1819), .b(n100), .O(n1820));
  nor2   g1756(.a(n1820), .b(n1818), .O(n1821));
  inv1   g1757(.a(n1821), .O(n1822));
  nor2   g1758(.a(n1822), .b(n1815), .O(n1823));
  inv1   g1759(.a(n1815), .O(n1824));
  nor2   g1760(.a(n1821), .b(n1824), .O(n1825));
  nor2   g1761(.a(n1825), .b(n1823), .O(n1826));
  inv1   g1762(.a(n1826), .O(n1827));
  nor2   g1763(.a(n1827), .b(n1814), .O(n1828));
  inv1   g1764(.a(n1814), .O(n1829));
  nor2   g1765(.a(n1826), .b(n1829), .O(n1830));
  nor2   g1766(.a(n1830), .b(n1828), .O(n1831));
  inv1   g1767(.a(n1831), .O(n1832));
  nor2   g1768(.a(n1832), .b(n1813), .O(n1833));
  inv1   g1769(.a(n1813), .O(n1834));
  nor2   g1770(.a(n1831), .b(n1834), .O(n1835));
  nor2   g1771(.a(n1835), .b(n1833), .O(n1836));
  inv1   g1772(.a(n1836), .O(n1837));
  nor2   g1773(.a(n1837), .b(n1812), .O(n1838));
  inv1   g1774(.a(n1812), .O(n1839));
  nor2   g1775(.a(n1836), .b(n1839), .O(n1840));
  nor2   g1776(.a(n1840), .b(n1838), .O(n1841));
  inv1   g1777(.a(n1841), .O(n1842));
  nor2   g1778(.a(n1842), .b(n1811), .O(n1843));
  inv1   g1779(.a(n1811), .O(n1844));
  nor2   g1780(.a(n1841), .b(n1844), .O(n1845));
  nor2   g1781(.a(n1845), .b(n1843), .O(n1846));
  inv1   g1782(.a(n1846), .O(n1847));
  nor2   g1783(.a(n1847), .b(n1810), .O(n1848));
  inv1   g1784(.a(n1810), .O(n1849));
  nor2   g1785(.a(n1846), .b(n1849), .O(n1850));
  nor2   g1786(.a(n1850), .b(n1848), .O(n1851));
  inv1   g1787(.a(n1851), .O(n1852));
  nor2   g1788(.a(n1852), .b(n1809), .O(n1853));
  inv1   g1789(.a(n1809), .O(n1854));
  nor2   g1790(.a(n1851), .b(n1854), .O(n1855));
  nor2   g1791(.a(n1855), .b(n1853), .O(n1856));
  inv1   g1792(.a(n1856), .O(n1857));
  nor2   g1793(.a(n1857), .b(n1808), .O(n1858));
  inv1   g1794(.a(n1808), .O(n1859));
  nor2   g1795(.a(n1856), .b(n1859), .O(n1860));
  nor2   g1796(.a(n1860), .b(n1858), .O(n1861));
  inv1   g1797(.a(n1861), .O(n1862));
  nor2   g1798(.a(n1862), .b(n1807), .O(n1863));
  inv1   g1799(.a(n1807), .O(n1864));
  nor2   g1800(.a(n1861), .b(n1864), .O(n1865));
  nor2   g1801(.a(n1865), .b(n1863), .O(n1866));
  inv1   g1802(.a(n1866), .O(n1867));
  nor2   g1803(.a(n1867), .b(n1806), .O(n1868));
  inv1   g1804(.a(n1806), .O(n1869));
  nor2   g1805(.a(n1866), .b(n1869), .O(n1870));
  nor2   g1806(.a(n1870), .b(n1868), .O(n1871));
  inv1   g1807(.a(n1871), .O(n1872));
  nor2   g1808(.a(n1872), .b(n1805), .O(n1873));
  inv1   g1809(.a(n1805), .O(n1874));
  nor2   g1810(.a(n1871), .b(n1874), .O(n1875));
  nor2   g1811(.a(n1875), .b(n1873), .O(n1876));
  inv1   g1812(.a(n1876), .O(n1877));
  nor2   g1813(.a(n1877), .b(n1804), .O(n1878));
  inv1   g1814(.a(n1804), .O(n1879));
  nor2   g1815(.a(n1876), .b(n1879), .O(n1880));
  nor2   g1816(.a(n1880), .b(n1878), .O(n1881));
  inv1   g1817(.a(n1881), .O(n1882));
  nor2   g1818(.a(n1882), .b(n1803), .O(n1883));
  inv1   g1819(.a(n1803), .O(n1884));
  nor2   g1820(.a(n1881), .b(n1884), .O(n1885));
  nor2   g1821(.a(n1885), .b(n1883), .O(n1886));
  inv1   g1822(.a(n1886), .O(n1887));
  nor2   g1823(.a(n1887), .b(n1802), .O(n1888));
  inv1   g1824(.a(n1802), .O(n1889));
  nor2   g1825(.a(n1886), .b(n1889), .O(n1890));
  nor2   g1826(.a(n1890), .b(n1888), .O(n1891));
  inv1   g1827(.a(n1891), .O(n1892));
  nor2   g1828(.a(n1892), .b(n1801), .O(n1893));
  inv1   g1829(.a(n1801), .O(n1894));
  nor2   g1830(.a(n1891), .b(n1894), .O(n1895));
  nor2   g1831(.a(n1895), .b(n1893), .O(n1896));
  inv1   g1832(.a(n1896), .O(n1897));
  nor2   g1833(.a(n1897), .b(n1800), .O(n1898));
  inv1   g1834(.a(n1800), .O(n1899));
  nor2   g1835(.a(n1896), .b(n1899), .O(n1900));
  nor2   g1836(.a(n1900), .b(n1898), .O(n1901));
  inv1   g1837(.a(n1901), .O(n1902));
  nor2   g1838(.a(n1902), .b(n1799), .O(n1903));
  inv1   g1839(.a(n1799), .O(n1904));
  nor2   g1840(.a(n1901), .b(n1904), .O(n1905));
  nor2   g1841(.a(n1905), .b(n1903), .O(n1906));
  inv1   g1842(.a(n1906), .O(n1907));
  nor2   g1843(.a(n1907), .b(n1798), .O(n1908));
  inv1   g1844(.a(n1798), .O(n1909));
  nor2   g1845(.a(n1906), .b(n1909), .O(n1910));
  nor2   g1846(.a(n1910), .b(n1908), .O(n1911));
  inv1   g1847(.a(n1911), .O(n1912));
  nor2   g1848(.a(n1912), .b(n1797), .O(n1913));
  inv1   g1849(.a(n1797), .O(n1914));
  nor2   g1850(.a(n1911), .b(n1914), .O(n1915));
  nor2   g1851(.a(n1915), .b(n1913), .O(n1916));
  inv1   g1852(.a(n1916), .O(n1917));
  nor2   g1853(.a(n1917), .b(n1796), .O(n1918));
  inv1   g1854(.a(n1796), .O(n1919));
  nor2   g1855(.a(n1916), .b(n1919), .O(n1920));
  nor2   g1856(.a(n1920), .b(n1918), .O(n1921));
  inv1   g1857(.a(n1921), .O(n1922));
  nor2   g1858(.a(n1922), .b(n1795), .O(n1923));
  inv1   g1859(.a(n1795), .O(n1924));
  nor2   g1860(.a(n1921), .b(n1924), .O(n1925));
  nor2   g1861(.a(n1925), .b(n1923), .O(n1926));
  inv1   g1862(.a(n1926), .O(n1927));
  nor2   g1863(.a(n1927), .b(n1794), .O(n1928));
  inv1   g1864(.a(n1794), .O(n1929));
  nor2   g1865(.a(n1926), .b(n1929), .O(n1930));
  nor2   g1866(.a(n1930), .b(n1928), .O(n1931));
  inv1   g1867(.a(n1931), .O(n1932));
  nor2   g1868(.a(n1932), .b(n1793), .O(n1933));
  inv1   g1869(.a(n1793), .O(n1934));
  nor2   g1870(.a(n1931), .b(n1934), .O(n1935));
  nor2   g1871(.a(n1935), .b(n1933), .O(n1936));
  inv1   g1872(.a(n1936), .O(n1937));
  nor2   g1873(.a(n1937), .b(n1792), .O(n1938));
  inv1   g1874(.a(n1792), .O(n1939));
  nor2   g1875(.a(n1936), .b(n1939), .O(n1940));
  nor2   g1876(.a(n1940), .b(n1938), .O(n1941));
  inv1   g1877(.a(n1941), .O(n1942));
  nor2   g1878(.a(n1942), .b(n1791), .O(n1943));
  inv1   g1879(.a(n1791), .O(n1944));
  nor2   g1880(.a(n1941), .b(n1944), .O(n1945));
  nor2   g1881(.a(n1945), .b(n1943), .O(n1946));
  inv1   g1882(.a(n1946), .O(G6170gat));
  nor2   g1883(.a(n1943), .b(n1938), .O(n1948));
  nor2   g1884(.a(n1933), .b(n1928), .O(n1949));
  nor2   g1885(.a(n1275), .b(n138), .O(n1950));
  nor2   g1886(.a(n1923), .b(n1918), .O(n1951));
  nor2   g1887(.a(n1111), .b(n184), .O(n1952));
  nor2   g1888(.a(n1913), .b(n1908), .O(n1953));
  nor2   g1889(.a(n959), .b(n242), .O(n1954));
  nor2   g1890(.a(n1903), .b(n1898), .O(n1955));
  nor2   g1891(.a(n819), .b(n312), .O(n1956));
  nor2   g1892(.a(n1893), .b(n1888), .O(n1957));
  nor2   g1893(.a(n691), .b(n394), .O(n1958));
  nor2   g1894(.a(n1883), .b(n1878), .O(n1959));
  nor2   g1895(.a(n575), .b(n488), .O(n1960));
  nor2   g1896(.a(n1873), .b(n1868), .O(n1961));
  nor2   g1897(.a(n471), .b(n594), .O(n1962));
  nor2   g1898(.a(n1863), .b(n1858), .O(n1963));
  nor2   g1899(.a(n379), .b(n712), .O(n1964));
  nor2   g1900(.a(n1853), .b(n1848), .O(n1965));
  nor2   g1901(.a(n299), .b(n842), .O(n1966));
  nor2   g1902(.a(n1843), .b(n1838), .O(n1967));
  nor2   g1903(.a(n231), .b(n984), .O(n1968));
  nor2   g1904(.a(n1833), .b(n1828), .O(n1969));
  nor2   g1905(.a(n175), .b(n1138), .O(n1970));
  nor2   g1906(.a(n131), .b(n1304), .O(n1971));
  nor2   g1907(.a(n1823), .b(n1818), .O(n1972));
  nor2   g1908(.a(n1972), .b(n1971), .O(n1973));
  inv1   g1909(.a(n1971), .O(n1974));
  inv1   g1910(.a(n1972), .O(n1975));
  nor2   g1911(.a(n1975), .b(n1974), .O(n1976));
  nor2   g1912(.a(n1976), .b(n1973), .O(n1977));
  inv1   g1913(.a(n1977), .O(n1978));
  nor2   g1914(.a(n1978), .b(n1970), .O(n1979));
  inv1   g1915(.a(n1970), .O(n1980));
  nor2   g1916(.a(n1977), .b(n1980), .O(n1981));
  nor2   g1917(.a(n1981), .b(n1979), .O(n1982));
  inv1   g1918(.a(n1982), .O(n1983));
  nor2   g1919(.a(n1983), .b(n1969), .O(n1984));
  inv1   g1920(.a(n1969), .O(n1985));
  nor2   g1921(.a(n1982), .b(n1985), .O(n1986));
  nor2   g1922(.a(n1986), .b(n1984), .O(n1987));
  inv1   g1923(.a(n1987), .O(n1988));
  nor2   g1924(.a(n1988), .b(n1968), .O(n1989));
  inv1   g1925(.a(n1968), .O(n1990));
  nor2   g1926(.a(n1987), .b(n1990), .O(n1991));
  nor2   g1927(.a(n1991), .b(n1989), .O(n1992));
  inv1   g1928(.a(n1992), .O(n1993));
  nor2   g1929(.a(n1993), .b(n1967), .O(n1994));
  inv1   g1930(.a(n1967), .O(n1995));
  nor2   g1931(.a(n1992), .b(n1995), .O(n1996));
  nor2   g1932(.a(n1996), .b(n1994), .O(n1997));
  inv1   g1933(.a(n1997), .O(n1998));
  nor2   g1934(.a(n1998), .b(n1966), .O(n1999));
  inv1   g1935(.a(n1966), .O(n2000));
  nor2   g1936(.a(n1997), .b(n2000), .O(n2001));
  nor2   g1937(.a(n2001), .b(n1999), .O(n2002));
  inv1   g1938(.a(n2002), .O(n2003));
  nor2   g1939(.a(n2003), .b(n1965), .O(n2004));
  inv1   g1940(.a(n1965), .O(n2005));
  nor2   g1941(.a(n2002), .b(n2005), .O(n2006));
  nor2   g1942(.a(n2006), .b(n2004), .O(n2007));
  inv1   g1943(.a(n2007), .O(n2008));
  nor2   g1944(.a(n2008), .b(n1964), .O(n2009));
  inv1   g1945(.a(n1964), .O(n2010));
  nor2   g1946(.a(n2007), .b(n2010), .O(n2011));
  nor2   g1947(.a(n2011), .b(n2009), .O(n2012));
  inv1   g1948(.a(n2012), .O(n2013));
  nor2   g1949(.a(n2013), .b(n1963), .O(n2014));
  inv1   g1950(.a(n1963), .O(n2015));
  nor2   g1951(.a(n2012), .b(n2015), .O(n2016));
  nor2   g1952(.a(n2016), .b(n2014), .O(n2017));
  inv1   g1953(.a(n2017), .O(n2018));
  nor2   g1954(.a(n2018), .b(n1962), .O(n2019));
  inv1   g1955(.a(n1962), .O(n2020));
  nor2   g1956(.a(n2017), .b(n2020), .O(n2021));
  nor2   g1957(.a(n2021), .b(n2019), .O(n2022));
  inv1   g1958(.a(n2022), .O(n2023));
  nor2   g1959(.a(n2023), .b(n1961), .O(n2024));
  inv1   g1960(.a(n1961), .O(n2025));
  nor2   g1961(.a(n2022), .b(n2025), .O(n2026));
  nor2   g1962(.a(n2026), .b(n2024), .O(n2027));
  inv1   g1963(.a(n2027), .O(n2028));
  nor2   g1964(.a(n2028), .b(n1960), .O(n2029));
  inv1   g1965(.a(n1960), .O(n2030));
  nor2   g1966(.a(n2027), .b(n2030), .O(n2031));
  nor2   g1967(.a(n2031), .b(n2029), .O(n2032));
  inv1   g1968(.a(n2032), .O(n2033));
  nor2   g1969(.a(n2033), .b(n1959), .O(n2034));
  inv1   g1970(.a(n1959), .O(n2035));
  nor2   g1971(.a(n2032), .b(n2035), .O(n2036));
  nor2   g1972(.a(n2036), .b(n2034), .O(n2037));
  inv1   g1973(.a(n2037), .O(n2038));
  nor2   g1974(.a(n2038), .b(n1958), .O(n2039));
  inv1   g1975(.a(n1958), .O(n2040));
  nor2   g1976(.a(n2037), .b(n2040), .O(n2041));
  nor2   g1977(.a(n2041), .b(n2039), .O(n2042));
  inv1   g1978(.a(n2042), .O(n2043));
  nor2   g1979(.a(n2043), .b(n1957), .O(n2044));
  inv1   g1980(.a(n1957), .O(n2045));
  nor2   g1981(.a(n2042), .b(n2045), .O(n2046));
  nor2   g1982(.a(n2046), .b(n2044), .O(n2047));
  inv1   g1983(.a(n2047), .O(n2048));
  nor2   g1984(.a(n2048), .b(n1956), .O(n2049));
  inv1   g1985(.a(n1956), .O(n2050));
  nor2   g1986(.a(n2047), .b(n2050), .O(n2051));
  nor2   g1987(.a(n2051), .b(n2049), .O(n2052));
  inv1   g1988(.a(n2052), .O(n2053));
  nor2   g1989(.a(n2053), .b(n1955), .O(n2054));
  inv1   g1990(.a(n1955), .O(n2055));
  nor2   g1991(.a(n2052), .b(n2055), .O(n2056));
  nor2   g1992(.a(n2056), .b(n2054), .O(n2057));
  inv1   g1993(.a(n2057), .O(n2058));
  nor2   g1994(.a(n2058), .b(n1954), .O(n2059));
  inv1   g1995(.a(n1954), .O(n2060));
  nor2   g1996(.a(n2057), .b(n2060), .O(n2061));
  nor2   g1997(.a(n2061), .b(n2059), .O(n2062));
  inv1   g1998(.a(n2062), .O(n2063));
  nor2   g1999(.a(n2063), .b(n1953), .O(n2064));
  inv1   g2000(.a(n1953), .O(n2065));
  nor2   g2001(.a(n2062), .b(n2065), .O(n2066));
  nor2   g2002(.a(n2066), .b(n2064), .O(n2067));
  inv1   g2003(.a(n2067), .O(n2068));
  nor2   g2004(.a(n2068), .b(n1952), .O(n2069));
  inv1   g2005(.a(n1952), .O(n2070));
  nor2   g2006(.a(n2067), .b(n2070), .O(n2071));
  nor2   g2007(.a(n2071), .b(n2069), .O(n2072));
  inv1   g2008(.a(n2072), .O(n2073));
  nor2   g2009(.a(n2073), .b(n1951), .O(n2074));
  inv1   g2010(.a(n1951), .O(n2075));
  nor2   g2011(.a(n2072), .b(n2075), .O(n2076));
  nor2   g2012(.a(n2076), .b(n2074), .O(n2077));
  inv1   g2013(.a(n2077), .O(n2078));
  nor2   g2014(.a(n2078), .b(n1950), .O(n2079));
  inv1   g2015(.a(n1950), .O(n2080));
  nor2   g2016(.a(n2077), .b(n2080), .O(n2081));
  nor2   g2017(.a(n2081), .b(n2079), .O(n2082));
  inv1   g2018(.a(n2082), .O(n2083));
  nor2   g2019(.a(n2083), .b(n1949), .O(n2084));
  inv1   g2020(.a(n1949), .O(n2085));
  nor2   g2021(.a(n2082), .b(n2085), .O(n2086));
  nor2   g2022(.a(n2086), .b(n2084), .O(n2087));
  inv1   g2023(.a(n2087), .O(n2088));
  nor2   g2024(.a(n2088), .b(n1948), .O(n2089));
  inv1   g2025(.a(n1948), .O(n2090));
  nor2   g2026(.a(n2087), .b(n2090), .O(n2091));
  nor2   g2027(.a(n2091), .b(n2089), .O(n2092));
  inv1   g2028(.a(n2092), .O(G6180gat));
  nor2   g2029(.a(n2089), .b(n2084), .O(n2094));
  nor2   g2030(.a(n2079), .b(n2074), .O(n2095));
  nor2   g2031(.a(n1275), .b(n184), .O(n2096));
  nor2   g2032(.a(n2069), .b(n2064), .O(n2097));
  nor2   g2033(.a(n1111), .b(n242), .O(n2098));
  nor2   g2034(.a(n2059), .b(n2054), .O(n2099));
  nor2   g2035(.a(n959), .b(n312), .O(n2100));
  nor2   g2036(.a(n2049), .b(n2044), .O(n2101));
  nor2   g2037(.a(n819), .b(n394), .O(n2102));
  nor2   g2038(.a(n2039), .b(n2034), .O(n2103));
  nor2   g2039(.a(n691), .b(n488), .O(n2104));
  nor2   g2040(.a(n2029), .b(n2024), .O(n2105));
  nor2   g2041(.a(n575), .b(n594), .O(n2106));
  nor2   g2042(.a(n2019), .b(n2014), .O(n2107));
  nor2   g2043(.a(n471), .b(n712), .O(n2108));
  nor2   g2044(.a(n2009), .b(n2004), .O(n2109));
  nor2   g2045(.a(n379), .b(n842), .O(n2110));
  nor2   g2046(.a(n1999), .b(n1994), .O(n2111));
  nor2   g2047(.a(n299), .b(n984), .O(n2112));
  nor2   g2048(.a(n1989), .b(n1984), .O(n2113));
  nor2   g2049(.a(n231), .b(n1138), .O(n2114));
  nor2   g2050(.a(n175), .b(n1304), .O(n2115));
  nor2   g2051(.a(n1979), .b(n1973), .O(n2116));
  nor2   g2052(.a(n2116), .b(n2115), .O(n2117));
  inv1   g2053(.a(n2115), .O(n2118));
  inv1   g2054(.a(n2116), .O(n2119));
  nor2   g2055(.a(n2119), .b(n2118), .O(n2120));
  nor2   g2056(.a(n2120), .b(n2117), .O(n2121));
  inv1   g2057(.a(n2121), .O(n2122));
  nor2   g2058(.a(n2122), .b(n2114), .O(n2123));
  inv1   g2059(.a(n2114), .O(n2124));
  nor2   g2060(.a(n2121), .b(n2124), .O(n2125));
  nor2   g2061(.a(n2125), .b(n2123), .O(n2126));
  inv1   g2062(.a(n2126), .O(n2127));
  nor2   g2063(.a(n2127), .b(n2113), .O(n2128));
  inv1   g2064(.a(n2113), .O(n2129));
  nor2   g2065(.a(n2126), .b(n2129), .O(n2130));
  nor2   g2066(.a(n2130), .b(n2128), .O(n2131));
  inv1   g2067(.a(n2131), .O(n2132));
  nor2   g2068(.a(n2132), .b(n2112), .O(n2133));
  inv1   g2069(.a(n2112), .O(n2134));
  nor2   g2070(.a(n2131), .b(n2134), .O(n2135));
  nor2   g2071(.a(n2135), .b(n2133), .O(n2136));
  inv1   g2072(.a(n2136), .O(n2137));
  nor2   g2073(.a(n2137), .b(n2111), .O(n2138));
  inv1   g2074(.a(n2111), .O(n2139));
  nor2   g2075(.a(n2136), .b(n2139), .O(n2140));
  nor2   g2076(.a(n2140), .b(n2138), .O(n2141));
  inv1   g2077(.a(n2141), .O(n2142));
  nor2   g2078(.a(n2142), .b(n2110), .O(n2143));
  inv1   g2079(.a(n2110), .O(n2144));
  nor2   g2080(.a(n2141), .b(n2144), .O(n2145));
  nor2   g2081(.a(n2145), .b(n2143), .O(n2146));
  inv1   g2082(.a(n2146), .O(n2147));
  nor2   g2083(.a(n2147), .b(n2109), .O(n2148));
  inv1   g2084(.a(n2109), .O(n2149));
  nor2   g2085(.a(n2146), .b(n2149), .O(n2150));
  nor2   g2086(.a(n2150), .b(n2148), .O(n2151));
  inv1   g2087(.a(n2151), .O(n2152));
  nor2   g2088(.a(n2152), .b(n2108), .O(n2153));
  inv1   g2089(.a(n2108), .O(n2154));
  nor2   g2090(.a(n2151), .b(n2154), .O(n2155));
  nor2   g2091(.a(n2155), .b(n2153), .O(n2156));
  inv1   g2092(.a(n2156), .O(n2157));
  nor2   g2093(.a(n2157), .b(n2107), .O(n2158));
  inv1   g2094(.a(n2107), .O(n2159));
  nor2   g2095(.a(n2156), .b(n2159), .O(n2160));
  nor2   g2096(.a(n2160), .b(n2158), .O(n2161));
  inv1   g2097(.a(n2161), .O(n2162));
  nor2   g2098(.a(n2162), .b(n2106), .O(n2163));
  inv1   g2099(.a(n2106), .O(n2164));
  nor2   g2100(.a(n2161), .b(n2164), .O(n2165));
  nor2   g2101(.a(n2165), .b(n2163), .O(n2166));
  inv1   g2102(.a(n2166), .O(n2167));
  nor2   g2103(.a(n2167), .b(n2105), .O(n2168));
  inv1   g2104(.a(n2105), .O(n2169));
  nor2   g2105(.a(n2166), .b(n2169), .O(n2170));
  nor2   g2106(.a(n2170), .b(n2168), .O(n2171));
  inv1   g2107(.a(n2171), .O(n2172));
  nor2   g2108(.a(n2172), .b(n2104), .O(n2173));
  inv1   g2109(.a(n2104), .O(n2174));
  nor2   g2110(.a(n2171), .b(n2174), .O(n2175));
  nor2   g2111(.a(n2175), .b(n2173), .O(n2176));
  inv1   g2112(.a(n2176), .O(n2177));
  nor2   g2113(.a(n2177), .b(n2103), .O(n2178));
  inv1   g2114(.a(n2103), .O(n2179));
  nor2   g2115(.a(n2176), .b(n2179), .O(n2180));
  nor2   g2116(.a(n2180), .b(n2178), .O(n2181));
  inv1   g2117(.a(n2181), .O(n2182));
  nor2   g2118(.a(n2182), .b(n2102), .O(n2183));
  inv1   g2119(.a(n2102), .O(n2184));
  nor2   g2120(.a(n2181), .b(n2184), .O(n2185));
  nor2   g2121(.a(n2185), .b(n2183), .O(n2186));
  inv1   g2122(.a(n2186), .O(n2187));
  nor2   g2123(.a(n2187), .b(n2101), .O(n2188));
  inv1   g2124(.a(n2101), .O(n2189));
  nor2   g2125(.a(n2186), .b(n2189), .O(n2190));
  nor2   g2126(.a(n2190), .b(n2188), .O(n2191));
  inv1   g2127(.a(n2191), .O(n2192));
  nor2   g2128(.a(n2192), .b(n2100), .O(n2193));
  inv1   g2129(.a(n2100), .O(n2194));
  nor2   g2130(.a(n2191), .b(n2194), .O(n2195));
  nor2   g2131(.a(n2195), .b(n2193), .O(n2196));
  inv1   g2132(.a(n2196), .O(n2197));
  nor2   g2133(.a(n2197), .b(n2099), .O(n2198));
  inv1   g2134(.a(n2099), .O(n2199));
  nor2   g2135(.a(n2196), .b(n2199), .O(n2200));
  nor2   g2136(.a(n2200), .b(n2198), .O(n2201));
  inv1   g2137(.a(n2201), .O(n2202));
  nor2   g2138(.a(n2202), .b(n2098), .O(n2203));
  inv1   g2139(.a(n2098), .O(n2204));
  nor2   g2140(.a(n2201), .b(n2204), .O(n2205));
  nor2   g2141(.a(n2205), .b(n2203), .O(n2206));
  inv1   g2142(.a(n2206), .O(n2207));
  nor2   g2143(.a(n2207), .b(n2097), .O(n2208));
  inv1   g2144(.a(n2097), .O(n2209));
  nor2   g2145(.a(n2206), .b(n2209), .O(n2210));
  nor2   g2146(.a(n2210), .b(n2208), .O(n2211));
  inv1   g2147(.a(n2211), .O(n2212));
  nor2   g2148(.a(n2212), .b(n2096), .O(n2213));
  inv1   g2149(.a(n2096), .O(n2214));
  nor2   g2150(.a(n2211), .b(n2214), .O(n2215));
  nor2   g2151(.a(n2215), .b(n2213), .O(n2216));
  inv1   g2152(.a(n2216), .O(n2217));
  nor2   g2153(.a(n2217), .b(n2095), .O(n2218));
  inv1   g2154(.a(n2095), .O(n2219));
  nor2   g2155(.a(n2216), .b(n2219), .O(n2220));
  nor2   g2156(.a(n2220), .b(n2218), .O(n2221));
  inv1   g2157(.a(n2221), .O(n2222));
  nor2   g2158(.a(n2222), .b(n2094), .O(n2223));
  inv1   g2159(.a(n2094), .O(n2224));
  nor2   g2160(.a(n2221), .b(n2224), .O(n2225));
  nor2   g2161(.a(n2225), .b(n2223), .O(n2226));
  inv1   g2162(.a(n2226), .O(G6190gat));
  nor2   g2163(.a(n2223), .b(n2218), .O(n2228));
  nor2   g2164(.a(n2213), .b(n2208), .O(n2229));
  nor2   g2165(.a(n1275), .b(n242), .O(n2230));
  nor2   g2166(.a(n2203), .b(n2198), .O(n2231));
  nor2   g2167(.a(n1111), .b(n312), .O(n2232));
  nor2   g2168(.a(n2193), .b(n2188), .O(n2233));
  nor2   g2169(.a(n959), .b(n394), .O(n2234));
  nor2   g2170(.a(n2183), .b(n2178), .O(n2235));
  nor2   g2171(.a(n819), .b(n488), .O(n2236));
  nor2   g2172(.a(n2173), .b(n2168), .O(n2237));
  nor2   g2173(.a(n691), .b(n594), .O(n2238));
  nor2   g2174(.a(n2163), .b(n2158), .O(n2239));
  nor2   g2175(.a(n575), .b(n712), .O(n2240));
  nor2   g2176(.a(n2153), .b(n2148), .O(n2241));
  nor2   g2177(.a(n471), .b(n842), .O(n2242));
  nor2   g2178(.a(n2143), .b(n2138), .O(n2243));
  nor2   g2179(.a(n379), .b(n984), .O(n2244));
  nor2   g2180(.a(n2133), .b(n2128), .O(n2245));
  nor2   g2181(.a(n299), .b(n1138), .O(n2246));
  nor2   g2182(.a(n231), .b(n1304), .O(n2247));
  nor2   g2183(.a(n2123), .b(n2117), .O(n2248));
  nor2   g2184(.a(n2248), .b(n2247), .O(n2249));
  inv1   g2185(.a(n2247), .O(n2250));
  inv1   g2186(.a(n2248), .O(n2251));
  nor2   g2187(.a(n2251), .b(n2250), .O(n2252));
  nor2   g2188(.a(n2252), .b(n2249), .O(n2253));
  inv1   g2189(.a(n2253), .O(n2254));
  nor2   g2190(.a(n2254), .b(n2246), .O(n2255));
  inv1   g2191(.a(n2246), .O(n2256));
  nor2   g2192(.a(n2253), .b(n2256), .O(n2257));
  nor2   g2193(.a(n2257), .b(n2255), .O(n2258));
  inv1   g2194(.a(n2258), .O(n2259));
  nor2   g2195(.a(n2259), .b(n2245), .O(n2260));
  inv1   g2196(.a(n2245), .O(n2261));
  nor2   g2197(.a(n2258), .b(n2261), .O(n2262));
  nor2   g2198(.a(n2262), .b(n2260), .O(n2263));
  inv1   g2199(.a(n2263), .O(n2264));
  nor2   g2200(.a(n2264), .b(n2244), .O(n2265));
  inv1   g2201(.a(n2244), .O(n2266));
  nor2   g2202(.a(n2263), .b(n2266), .O(n2267));
  nor2   g2203(.a(n2267), .b(n2265), .O(n2268));
  inv1   g2204(.a(n2268), .O(n2269));
  nor2   g2205(.a(n2269), .b(n2243), .O(n2270));
  inv1   g2206(.a(n2243), .O(n2271));
  nor2   g2207(.a(n2268), .b(n2271), .O(n2272));
  nor2   g2208(.a(n2272), .b(n2270), .O(n2273));
  inv1   g2209(.a(n2273), .O(n2274));
  nor2   g2210(.a(n2274), .b(n2242), .O(n2275));
  inv1   g2211(.a(n2242), .O(n2276));
  nor2   g2212(.a(n2273), .b(n2276), .O(n2277));
  nor2   g2213(.a(n2277), .b(n2275), .O(n2278));
  inv1   g2214(.a(n2278), .O(n2279));
  nor2   g2215(.a(n2279), .b(n2241), .O(n2280));
  inv1   g2216(.a(n2241), .O(n2281));
  nor2   g2217(.a(n2278), .b(n2281), .O(n2282));
  nor2   g2218(.a(n2282), .b(n2280), .O(n2283));
  inv1   g2219(.a(n2283), .O(n2284));
  nor2   g2220(.a(n2284), .b(n2240), .O(n2285));
  inv1   g2221(.a(n2240), .O(n2286));
  nor2   g2222(.a(n2283), .b(n2286), .O(n2287));
  nor2   g2223(.a(n2287), .b(n2285), .O(n2288));
  inv1   g2224(.a(n2288), .O(n2289));
  nor2   g2225(.a(n2289), .b(n2239), .O(n2290));
  inv1   g2226(.a(n2239), .O(n2291));
  nor2   g2227(.a(n2288), .b(n2291), .O(n2292));
  nor2   g2228(.a(n2292), .b(n2290), .O(n2293));
  inv1   g2229(.a(n2293), .O(n2294));
  nor2   g2230(.a(n2294), .b(n2238), .O(n2295));
  inv1   g2231(.a(n2238), .O(n2296));
  nor2   g2232(.a(n2293), .b(n2296), .O(n2297));
  nor2   g2233(.a(n2297), .b(n2295), .O(n2298));
  inv1   g2234(.a(n2298), .O(n2299));
  nor2   g2235(.a(n2299), .b(n2237), .O(n2300));
  inv1   g2236(.a(n2237), .O(n2301));
  nor2   g2237(.a(n2298), .b(n2301), .O(n2302));
  nor2   g2238(.a(n2302), .b(n2300), .O(n2303));
  inv1   g2239(.a(n2303), .O(n2304));
  nor2   g2240(.a(n2304), .b(n2236), .O(n2305));
  inv1   g2241(.a(n2236), .O(n2306));
  nor2   g2242(.a(n2303), .b(n2306), .O(n2307));
  nor2   g2243(.a(n2307), .b(n2305), .O(n2308));
  inv1   g2244(.a(n2308), .O(n2309));
  nor2   g2245(.a(n2309), .b(n2235), .O(n2310));
  inv1   g2246(.a(n2235), .O(n2311));
  nor2   g2247(.a(n2308), .b(n2311), .O(n2312));
  nor2   g2248(.a(n2312), .b(n2310), .O(n2313));
  inv1   g2249(.a(n2313), .O(n2314));
  nor2   g2250(.a(n2314), .b(n2234), .O(n2315));
  inv1   g2251(.a(n2234), .O(n2316));
  nor2   g2252(.a(n2313), .b(n2316), .O(n2317));
  nor2   g2253(.a(n2317), .b(n2315), .O(n2318));
  inv1   g2254(.a(n2318), .O(n2319));
  nor2   g2255(.a(n2319), .b(n2233), .O(n2320));
  inv1   g2256(.a(n2233), .O(n2321));
  nor2   g2257(.a(n2318), .b(n2321), .O(n2322));
  nor2   g2258(.a(n2322), .b(n2320), .O(n2323));
  inv1   g2259(.a(n2323), .O(n2324));
  nor2   g2260(.a(n2324), .b(n2232), .O(n2325));
  inv1   g2261(.a(n2232), .O(n2326));
  nor2   g2262(.a(n2323), .b(n2326), .O(n2327));
  nor2   g2263(.a(n2327), .b(n2325), .O(n2328));
  inv1   g2264(.a(n2328), .O(n2329));
  nor2   g2265(.a(n2329), .b(n2231), .O(n2330));
  inv1   g2266(.a(n2231), .O(n2331));
  nor2   g2267(.a(n2328), .b(n2331), .O(n2332));
  nor2   g2268(.a(n2332), .b(n2330), .O(n2333));
  inv1   g2269(.a(n2333), .O(n2334));
  nor2   g2270(.a(n2334), .b(n2230), .O(n2335));
  inv1   g2271(.a(n2230), .O(n2336));
  nor2   g2272(.a(n2333), .b(n2336), .O(n2337));
  nor2   g2273(.a(n2337), .b(n2335), .O(n2338));
  inv1   g2274(.a(n2338), .O(n2339));
  nor2   g2275(.a(n2339), .b(n2229), .O(n2340));
  inv1   g2276(.a(n2229), .O(n2341));
  nor2   g2277(.a(n2338), .b(n2341), .O(n2342));
  nor2   g2278(.a(n2342), .b(n2340), .O(n2343));
  inv1   g2279(.a(n2343), .O(n2344));
  nor2   g2280(.a(n2344), .b(n2228), .O(n2345));
  inv1   g2281(.a(n2228), .O(n2346));
  nor2   g2282(.a(n2343), .b(n2346), .O(n2347));
  nor2   g2283(.a(n2347), .b(n2345), .O(n2348));
  inv1   g2284(.a(n2348), .O(G6200gat));
  nor2   g2285(.a(n2345), .b(n2340), .O(n2350));
  nor2   g2286(.a(n2335), .b(n2330), .O(n2351));
  nor2   g2287(.a(n1275), .b(n312), .O(n2352));
  nor2   g2288(.a(n2325), .b(n2320), .O(n2353));
  nor2   g2289(.a(n1111), .b(n394), .O(n2354));
  nor2   g2290(.a(n2315), .b(n2310), .O(n2355));
  nor2   g2291(.a(n959), .b(n488), .O(n2356));
  nor2   g2292(.a(n2305), .b(n2300), .O(n2357));
  nor2   g2293(.a(n819), .b(n594), .O(n2358));
  nor2   g2294(.a(n2295), .b(n2290), .O(n2359));
  nor2   g2295(.a(n691), .b(n712), .O(n2360));
  nor2   g2296(.a(n2285), .b(n2280), .O(n2361));
  nor2   g2297(.a(n575), .b(n842), .O(n2362));
  nor2   g2298(.a(n2275), .b(n2270), .O(n2363));
  nor2   g2299(.a(n471), .b(n984), .O(n2364));
  nor2   g2300(.a(n2265), .b(n2260), .O(n2365));
  nor2   g2301(.a(n379), .b(n1138), .O(n2366));
  nor2   g2302(.a(n299), .b(n1304), .O(n2367));
  nor2   g2303(.a(n2255), .b(n2249), .O(n2368));
  nor2   g2304(.a(n2368), .b(n2367), .O(n2369));
  inv1   g2305(.a(n2367), .O(n2370));
  inv1   g2306(.a(n2368), .O(n2371));
  nor2   g2307(.a(n2371), .b(n2370), .O(n2372));
  nor2   g2308(.a(n2372), .b(n2369), .O(n2373));
  inv1   g2309(.a(n2373), .O(n2374));
  nor2   g2310(.a(n2374), .b(n2366), .O(n2375));
  inv1   g2311(.a(n2366), .O(n2376));
  nor2   g2312(.a(n2373), .b(n2376), .O(n2377));
  nor2   g2313(.a(n2377), .b(n2375), .O(n2378));
  inv1   g2314(.a(n2378), .O(n2379));
  nor2   g2315(.a(n2379), .b(n2365), .O(n2380));
  inv1   g2316(.a(n2365), .O(n2381));
  nor2   g2317(.a(n2378), .b(n2381), .O(n2382));
  nor2   g2318(.a(n2382), .b(n2380), .O(n2383));
  inv1   g2319(.a(n2383), .O(n2384));
  nor2   g2320(.a(n2384), .b(n2364), .O(n2385));
  inv1   g2321(.a(n2364), .O(n2386));
  nor2   g2322(.a(n2383), .b(n2386), .O(n2387));
  nor2   g2323(.a(n2387), .b(n2385), .O(n2388));
  inv1   g2324(.a(n2388), .O(n2389));
  nor2   g2325(.a(n2389), .b(n2363), .O(n2390));
  inv1   g2326(.a(n2363), .O(n2391));
  nor2   g2327(.a(n2388), .b(n2391), .O(n2392));
  nor2   g2328(.a(n2392), .b(n2390), .O(n2393));
  inv1   g2329(.a(n2393), .O(n2394));
  nor2   g2330(.a(n2394), .b(n2362), .O(n2395));
  inv1   g2331(.a(n2362), .O(n2396));
  nor2   g2332(.a(n2393), .b(n2396), .O(n2397));
  nor2   g2333(.a(n2397), .b(n2395), .O(n2398));
  inv1   g2334(.a(n2398), .O(n2399));
  nor2   g2335(.a(n2399), .b(n2361), .O(n2400));
  inv1   g2336(.a(n2361), .O(n2401));
  nor2   g2337(.a(n2398), .b(n2401), .O(n2402));
  nor2   g2338(.a(n2402), .b(n2400), .O(n2403));
  inv1   g2339(.a(n2403), .O(n2404));
  nor2   g2340(.a(n2404), .b(n2360), .O(n2405));
  inv1   g2341(.a(n2360), .O(n2406));
  nor2   g2342(.a(n2403), .b(n2406), .O(n2407));
  nor2   g2343(.a(n2407), .b(n2405), .O(n2408));
  inv1   g2344(.a(n2408), .O(n2409));
  nor2   g2345(.a(n2409), .b(n2359), .O(n2410));
  inv1   g2346(.a(n2359), .O(n2411));
  nor2   g2347(.a(n2408), .b(n2411), .O(n2412));
  nor2   g2348(.a(n2412), .b(n2410), .O(n2413));
  inv1   g2349(.a(n2413), .O(n2414));
  nor2   g2350(.a(n2414), .b(n2358), .O(n2415));
  inv1   g2351(.a(n2358), .O(n2416));
  nor2   g2352(.a(n2413), .b(n2416), .O(n2417));
  nor2   g2353(.a(n2417), .b(n2415), .O(n2418));
  inv1   g2354(.a(n2418), .O(n2419));
  nor2   g2355(.a(n2419), .b(n2357), .O(n2420));
  inv1   g2356(.a(n2357), .O(n2421));
  nor2   g2357(.a(n2418), .b(n2421), .O(n2422));
  nor2   g2358(.a(n2422), .b(n2420), .O(n2423));
  inv1   g2359(.a(n2423), .O(n2424));
  nor2   g2360(.a(n2424), .b(n2356), .O(n2425));
  inv1   g2361(.a(n2356), .O(n2426));
  nor2   g2362(.a(n2423), .b(n2426), .O(n2427));
  nor2   g2363(.a(n2427), .b(n2425), .O(n2428));
  inv1   g2364(.a(n2428), .O(n2429));
  nor2   g2365(.a(n2429), .b(n2355), .O(n2430));
  inv1   g2366(.a(n2355), .O(n2431));
  nor2   g2367(.a(n2428), .b(n2431), .O(n2432));
  nor2   g2368(.a(n2432), .b(n2430), .O(n2433));
  inv1   g2369(.a(n2433), .O(n2434));
  nor2   g2370(.a(n2434), .b(n2354), .O(n2435));
  inv1   g2371(.a(n2354), .O(n2436));
  nor2   g2372(.a(n2433), .b(n2436), .O(n2437));
  nor2   g2373(.a(n2437), .b(n2435), .O(n2438));
  inv1   g2374(.a(n2438), .O(n2439));
  nor2   g2375(.a(n2439), .b(n2353), .O(n2440));
  inv1   g2376(.a(n2353), .O(n2441));
  nor2   g2377(.a(n2438), .b(n2441), .O(n2442));
  nor2   g2378(.a(n2442), .b(n2440), .O(n2443));
  inv1   g2379(.a(n2443), .O(n2444));
  nor2   g2380(.a(n2444), .b(n2352), .O(n2445));
  inv1   g2381(.a(n2352), .O(n2446));
  nor2   g2382(.a(n2443), .b(n2446), .O(n2447));
  nor2   g2383(.a(n2447), .b(n2445), .O(n2448));
  inv1   g2384(.a(n2448), .O(n2449));
  nor2   g2385(.a(n2449), .b(n2351), .O(n2450));
  inv1   g2386(.a(n2351), .O(n2451));
  nor2   g2387(.a(n2448), .b(n2451), .O(n2452));
  nor2   g2388(.a(n2452), .b(n2450), .O(n2453));
  inv1   g2389(.a(n2453), .O(n2454));
  nor2   g2390(.a(n2454), .b(n2350), .O(n2455));
  inv1   g2391(.a(n2350), .O(n2456));
  nor2   g2392(.a(n2453), .b(n2456), .O(n2457));
  nor2   g2393(.a(n2457), .b(n2455), .O(n2458));
  inv1   g2394(.a(n2458), .O(G6210gat));
  nor2   g2395(.a(n2455), .b(n2450), .O(n2460));
  nor2   g2396(.a(n2445), .b(n2440), .O(n2461));
  nor2   g2397(.a(n1275), .b(n394), .O(n2462));
  nor2   g2398(.a(n2435), .b(n2430), .O(n2463));
  nor2   g2399(.a(n1111), .b(n488), .O(n2464));
  nor2   g2400(.a(n2425), .b(n2420), .O(n2465));
  nor2   g2401(.a(n959), .b(n594), .O(n2466));
  nor2   g2402(.a(n2415), .b(n2410), .O(n2467));
  nor2   g2403(.a(n819), .b(n712), .O(n2468));
  nor2   g2404(.a(n2405), .b(n2400), .O(n2469));
  nor2   g2405(.a(n691), .b(n842), .O(n2470));
  nor2   g2406(.a(n2395), .b(n2390), .O(n2471));
  nor2   g2407(.a(n575), .b(n984), .O(n2472));
  nor2   g2408(.a(n2385), .b(n2380), .O(n2473));
  nor2   g2409(.a(n471), .b(n1138), .O(n2474));
  nor2   g2410(.a(n379), .b(n1304), .O(n2475));
  nor2   g2411(.a(n2375), .b(n2369), .O(n2476));
  nor2   g2412(.a(n2476), .b(n2475), .O(n2477));
  inv1   g2413(.a(n2475), .O(n2478));
  inv1   g2414(.a(n2476), .O(n2479));
  nor2   g2415(.a(n2479), .b(n2478), .O(n2480));
  nor2   g2416(.a(n2480), .b(n2477), .O(n2481));
  inv1   g2417(.a(n2481), .O(n2482));
  nor2   g2418(.a(n2482), .b(n2474), .O(n2483));
  inv1   g2419(.a(n2474), .O(n2484));
  nor2   g2420(.a(n2481), .b(n2484), .O(n2485));
  nor2   g2421(.a(n2485), .b(n2483), .O(n2486));
  inv1   g2422(.a(n2486), .O(n2487));
  nor2   g2423(.a(n2487), .b(n2473), .O(n2488));
  inv1   g2424(.a(n2473), .O(n2489));
  nor2   g2425(.a(n2486), .b(n2489), .O(n2490));
  nor2   g2426(.a(n2490), .b(n2488), .O(n2491));
  inv1   g2427(.a(n2491), .O(n2492));
  nor2   g2428(.a(n2492), .b(n2472), .O(n2493));
  inv1   g2429(.a(n2472), .O(n2494));
  nor2   g2430(.a(n2491), .b(n2494), .O(n2495));
  nor2   g2431(.a(n2495), .b(n2493), .O(n2496));
  inv1   g2432(.a(n2496), .O(n2497));
  nor2   g2433(.a(n2497), .b(n2471), .O(n2498));
  inv1   g2434(.a(n2471), .O(n2499));
  nor2   g2435(.a(n2496), .b(n2499), .O(n2500));
  nor2   g2436(.a(n2500), .b(n2498), .O(n2501));
  inv1   g2437(.a(n2501), .O(n2502));
  nor2   g2438(.a(n2502), .b(n2470), .O(n2503));
  inv1   g2439(.a(n2470), .O(n2504));
  nor2   g2440(.a(n2501), .b(n2504), .O(n2505));
  nor2   g2441(.a(n2505), .b(n2503), .O(n2506));
  inv1   g2442(.a(n2506), .O(n2507));
  nor2   g2443(.a(n2507), .b(n2469), .O(n2508));
  inv1   g2444(.a(n2469), .O(n2509));
  nor2   g2445(.a(n2506), .b(n2509), .O(n2510));
  nor2   g2446(.a(n2510), .b(n2508), .O(n2511));
  inv1   g2447(.a(n2511), .O(n2512));
  nor2   g2448(.a(n2512), .b(n2468), .O(n2513));
  inv1   g2449(.a(n2468), .O(n2514));
  nor2   g2450(.a(n2511), .b(n2514), .O(n2515));
  nor2   g2451(.a(n2515), .b(n2513), .O(n2516));
  inv1   g2452(.a(n2516), .O(n2517));
  nor2   g2453(.a(n2517), .b(n2467), .O(n2518));
  inv1   g2454(.a(n2467), .O(n2519));
  nor2   g2455(.a(n2516), .b(n2519), .O(n2520));
  nor2   g2456(.a(n2520), .b(n2518), .O(n2521));
  inv1   g2457(.a(n2521), .O(n2522));
  nor2   g2458(.a(n2522), .b(n2466), .O(n2523));
  inv1   g2459(.a(n2466), .O(n2524));
  nor2   g2460(.a(n2521), .b(n2524), .O(n2525));
  nor2   g2461(.a(n2525), .b(n2523), .O(n2526));
  inv1   g2462(.a(n2526), .O(n2527));
  nor2   g2463(.a(n2527), .b(n2465), .O(n2528));
  inv1   g2464(.a(n2465), .O(n2529));
  nor2   g2465(.a(n2526), .b(n2529), .O(n2530));
  nor2   g2466(.a(n2530), .b(n2528), .O(n2531));
  inv1   g2467(.a(n2531), .O(n2532));
  nor2   g2468(.a(n2532), .b(n2464), .O(n2533));
  inv1   g2469(.a(n2464), .O(n2534));
  nor2   g2470(.a(n2531), .b(n2534), .O(n2535));
  nor2   g2471(.a(n2535), .b(n2533), .O(n2536));
  inv1   g2472(.a(n2536), .O(n2537));
  nor2   g2473(.a(n2537), .b(n2463), .O(n2538));
  inv1   g2474(.a(n2463), .O(n2539));
  nor2   g2475(.a(n2536), .b(n2539), .O(n2540));
  nor2   g2476(.a(n2540), .b(n2538), .O(n2541));
  inv1   g2477(.a(n2541), .O(n2542));
  nor2   g2478(.a(n2542), .b(n2462), .O(n2543));
  inv1   g2479(.a(n2462), .O(n2544));
  nor2   g2480(.a(n2541), .b(n2544), .O(n2545));
  nor2   g2481(.a(n2545), .b(n2543), .O(n2546));
  inv1   g2482(.a(n2546), .O(n2547));
  nor2   g2483(.a(n2547), .b(n2461), .O(n2548));
  inv1   g2484(.a(n2461), .O(n2549));
  nor2   g2485(.a(n2546), .b(n2549), .O(n2550));
  nor2   g2486(.a(n2550), .b(n2548), .O(n2551));
  inv1   g2487(.a(n2551), .O(n2552));
  nor2   g2488(.a(n2552), .b(n2460), .O(n2553));
  inv1   g2489(.a(n2460), .O(n2554));
  nor2   g2490(.a(n2551), .b(n2554), .O(n2555));
  nor2   g2491(.a(n2555), .b(n2553), .O(n2556));
  inv1   g2492(.a(n2556), .O(G6220gat));
  nor2   g2493(.a(n2553), .b(n2548), .O(n2558));
  nor2   g2494(.a(n2543), .b(n2538), .O(n2559));
  nor2   g2495(.a(n1275), .b(n488), .O(n2560));
  nor2   g2496(.a(n2533), .b(n2528), .O(n2561));
  nor2   g2497(.a(n1111), .b(n594), .O(n2562));
  nor2   g2498(.a(n2523), .b(n2518), .O(n2563));
  nor2   g2499(.a(n959), .b(n712), .O(n2564));
  nor2   g2500(.a(n2513), .b(n2508), .O(n2565));
  nor2   g2501(.a(n819), .b(n842), .O(n2566));
  nor2   g2502(.a(n2503), .b(n2498), .O(n2567));
  nor2   g2503(.a(n691), .b(n984), .O(n2568));
  nor2   g2504(.a(n2493), .b(n2488), .O(n2569));
  nor2   g2505(.a(n575), .b(n1138), .O(n2570));
  nor2   g2506(.a(n471), .b(n1304), .O(n2571));
  nor2   g2507(.a(n2483), .b(n2477), .O(n2572));
  nor2   g2508(.a(n2572), .b(n2571), .O(n2573));
  inv1   g2509(.a(n2571), .O(n2574));
  inv1   g2510(.a(n2572), .O(n2575));
  nor2   g2511(.a(n2575), .b(n2574), .O(n2576));
  nor2   g2512(.a(n2576), .b(n2573), .O(n2577));
  inv1   g2513(.a(n2577), .O(n2578));
  nor2   g2514(.a(n2578), .b(n2570), .O(n2579));
  inv1   g2515(.a(n2570), .O(n2580));
  nor2   g2516(.a(n2577), .b(n2580), .O(n2581));
  nor2   g2517(.a(n2581), .b(n2579), .O(n2582));
  inv1   g2518(.a(n2582), .O(n2583));
  nor2   g2519(.a(n2583), .b(n2569), .O(n2584));
  inv1   g2520(.a(n2569), .O(n2585));
  nor2   g2521(.a(n2582), .b(n2585), .O(n2586));
  nor2   g2522(.a(n2586), .b(n2584), .O(n2587));
  inv1   g2523(.a(n2587), .O(n2588));
  nor2   g2524(.a(n2588), .b(n2568), .O(n2589));
  inv1   g2525(.a(n2568), .O(n2590));
  nor2   g2526(.a(n2587), .b(n2590), .O(n2591));
  nor2   g2527(.a(n2591), .b(n2589), .O(n2592));
  inv1   g2528(.a(n2592), .O(n2593));
  nor2   g2529(.a(n2593), .b(n2567), .O(n2594));
  inv1   g2530(.a(n2567), .O(n2595));
  nor2   g2531(.a(n2592), .b(n2595), .O(n2596));
  nor2   g2532(.a(n2596), .b(n2594), .O(n2597));
  inv1   g2533(.a(n2597), .O(n2598));
  nor2   g2534(.a(n2598), .b(n2566), .O(n2599));
  inv1   g2535(.a(n2566), .O(n2600));
  nor2   g2536(.a(n2597), .b(n2600), .O(n2601));
  nor2   g2537(.a(n2601), .b(n2599), .O(n2602));
  inv1   g2538(.a(n2602), .O(n2603));
  nor2   g2539(.a(n2603), .b(n2565), .O(n2604));
  inv1   g2540(.a(n2565), .O(n2605));
  nor2   g2541(.a(n2602), .b(n2605), .O(n2606));
  nor2   g2542(.a(n2606), .b(n2604), .O(n2607));
  inv1   g2543(.a(n2607), .O(n2608));
  nor2   g2544(.a(n2608), .b(n2564), .O(n2609));
  inv1   g2545(.a(n2564), .O(n2610));
  nor2   g2546(.a(n2607), .b(n2610), .O(n2611));
  nor2   g2547(.a(n2611), .b(n2609), .O(n2612));
  inv1   g2548(.a(n2612), .O(n2613));
  nor2   g2549(.a(n2613), .b(n2563), .O(n2614));
  inv1   g2550(.a(n2563), .O(n2615));
  nor2   g2551(.a(n2612), .b(n2615), .O(n2616));
  nor2   g2552(.a(n2616), .b(n2614), .O(n2617));
  inv1   g2553(.a(n2617), .O(n2618));
  nor2   g2554(.a(n2618), .b(n2562), .O(n2619));
  inv1   g2555(.a(n2562), .O(n2620));
  nor2   g2556(.a(n2617), .b(n2620), .O(n2621));
  nor2   g2557(.a(n2621), .b(n2619), .O(n2622));
  inv1   g2558(.a(n2622), .O(n2623));
  nor2   g2559(.a(n2623), .b(n2561), .O(n2624));
  inv1   g2560(.a(n2561), .O(n2625));
  nor2   g2561(.a(n2622), .b(n2625), .O(n2626));
  nor2   g2562(.a(n2626), .b(n2624), .O(n2627));
  inv1   g2563(.a(n2627), .O(n2628));
  nor2   g2564(.a(n2628), .b(n2560), .O(n2629));
  inv1   g2565(.a(n2560), .O(n2630));
  nor2   g2566(.a(n2627), .b(n2630), .O(n2631));
  nor2   g2567(.a(n2631), .b(n2629), .O(n2632));
  inv1   g2568(.a(n2632), .O(n2633));
  nor2   g2569(.a(n2633), .b(n2559), .O(n2634));
  inv1   g2570(.a(n2559), .O(n2635));
  nor2   g2571(.a(n2632), .b(n2635), .O(n2636));
  nor2   g2572(.a(n2636), .b(n2634), .O(n2637));
  inv1   g2573(.a(n2637), .O(n2638));
  nor2   g2574(.a(n2638), .b(n2558), .O(n2639));
  inv1   g2575(.a(n2558), .O(n2640));
  nor2   g2576(.a(n2637), .b(n2640), .O(n2641));
  nor2   g2577(.a(n2641), .b(n2639), .O(n2642));
  inv1   g2578(.a(n2642), .O(G6230gat));
  nor2   g2579(.a(n2639), .b(n2634), .O(n2644));
  nor2   g2580(.a(n2629), .b(n2624), .O(n2645));
  nor2   g2581(.a(n1275), .b(n594), .O(n2646));
  nor2   g2582(.a(n2619), .b(n2614), .O(n2647));
  nor2   g2583(.a(n1111), .b(n712), .O(n2648));
  nor2   g2584(.a(n2609), .b(n2604), .O(n2649));
  nor2   g2585(.a(n959), .b(n842), .O(n2650));
  nor2   g2586(.a(n2599), .b(n2594), .O(n2651));
  nor2   g2587(.a(n819), .b(n984), .O(n2652));
  nor2   g2588(.a(n2589), .b(n2584), .O(n2653));
  nor2   g2589(.a(n691), .b(n1138), .O(n2654));
  nor2   g2590(.a(n575), .b(n1304), .O(n2655));
  nor2   g2591(.a(n2579), .b(n2573), .O(n2656));
  nor2   g2592(.a(n2656), .b(n2655), .O(n2657));
  inv1   g2593(.a(n2655), .O(n2658));
  inv1   g2594(.a(n2656), .O(n2659));
  nor2   g2595(.a(n2659), .b(n2658), .O(n2660));
  nor2   g2596(.a(n2660), .b(n2657), .O(n2661));
  inv1   g2597(.a(n2661), .O(n2662));
  nor2   g2598(.a(n2662), .b(n2654), .O(n2663));
  inv1   g2599(.a(n2654), .O(n2664));
  nor2   g2600(.a(n2661), .b(n2664), .O(n2665));
  nor2   g2601(.a(n2665), .b(n2663), .O(n2666));
  inv1   g2602(.a(n2666), .O(n2667));
  nor2   g2603(.a(n2667), .b(n2653), .O(n2668));
  inv1   g2604(.a(n2653), .O(n2669));
  nor2   g2605(.a(n2666), .b(n2669), .O(n2670));
  nor2   g2606(.a(n2670), .b(n2668), .O(n2671));
  inv1   g2607(.a(n2671), .O(n2672));
  nor2   g2608(.a(n2672), .b(n2652), .O(n2673));
  inv1   g2609(.a(n2652), .O(n2674));
  nor2   g2610(.a(n2671), .b(n2674), .O(n2675));
  nor2   g2611(.a(n2675), .b(n2673), .O(n2676));
  inv1   g2612(.a(n2676), .O(n2677));
  nor2   g2613(.a(n2677), .b(n2651), .O(n2678));
  inv1   g2614(.a(n2651), .O(n2679));
  nor2   g2615(.a(n2676), .b(n2679), .O(n2680));
  nor2   g2616(.a(n2680), .b(n2678), .O(n2681));
  inv1   g2617(.a(n2681), .O(n2682));
  nor2   g2618(.a(n2682), .b(n2650), .O(n2683));
  inv1   g2619(.a(n2650), .O(n2684));
  nor2   g2620(.a(n2681), .b(n2684), .O(n2685));
  nor2   g2621(.a(n2685), .b(n2683), .O(n2686));
  inv1   g2622(.a(n2686), .O(n2687));
  nor2   g2623(.a(n2687), .b(n2649), .O(n2688));
  inv1   g2624(.a(n2649), .O(n2689));
  nor2   g2625(.a(n2686), .b(n2689), .O(n2690));
  nor2   g2626(.a(n2690), .b(n2688), .O(n2691));
  inv1   g2627(.a(n2691), .O(n2692));
  nor2   g2628(.a(n2692), .b(n2648), .O(n2693));
  inv1   g2629(.a(n2648), .O(n2694));
  nor2   g2630(.a(n2691), .b(n2694), .O(n2695));
  nor2   g2631(.a(n2695), .b(n2693), .O(n2696));
  inv1   g2632(.a(n2696), .O(n2697));
  nor2   g2633(.a(n2697), .b(n2647), .O(n2698));
  inv1   g2634(.a(n2647), .O(n2699));
  nor2   g2635(.a(n2696), .b(n2699), .O(n2700));
  nor2   g2636(.a(n2700), .b(n2698), .O(n2701));
  inv1   g2637(.a(n2701), .O(n2702));
  nor2   g2638(.a(n2702), .b(n2646), .O(n2703));
  inv1   g2639(.a(n2646), .O(n2704));
  nor2   g2640(.a(n2701), .b(n2704), .O(n2705));
  nor2   g2641(.a(n2705), .b(n2703), .O(n2706));
  inv1   g2642(.a(n2706), .O(n2707));
  nor2   g2643(.a(n2707), .b(n2645), .O(n2708));
  inv1   g2644(.a(n2645), .O(n2709));
  nor2   g2645(.a(n2706), .b(n2709), .O(n2710));
  nor2   g2646(.a(n2710), .b(n2708), .O(n2711));
  inv1   g2647(.a(n2711), .O(n2712));
  nor2   g2648(.a(n2712), .b(n2644), .O(n2713));
  inv1   g2649(.a(n2644), .O(n2714));
  nor2   g2650(.a(n2711), .b(n2714), .O(n2715));
  nor2   g2651(.a(n2715), .b(n2713), .O(n2716));
  inv1   g2652(.a(n2716), .O(G6240gat));
  nor2   g2653(.a(n2713), .b(n2708), .O(n2718));
  nor2   g2654(.a(n2703), .b(n2698), .O(n2719));
  nor2   g2655(.a(n1275), .b(n712), .O(n2720));
  nor2   g2656(.a(n2693), .b(n2688), .O(n2721));
  nor2   g2657(.a(n1111), .b(n842), .O(n2722));
  nor2   g2658(.a(n2683), .b(n2678), .O(n2723));
  nor2   g2659(.a(n959), .b(n984), .O(n2724));
  nor2   g2660(.a(n2673), .b(n2668), .O(n2725));
  nor2   g2661(.a(n819), .b(n1138), .O(n2726));
  nor2   g2662(.a(n691), .b(n1304), .O(n2727));
  nor2   g2663(.a(n2663), .b(n2657), .O(n2728));
  nor2   g2664(.a(n2728), .b(n2727), .O(n2729));
  inv1   g2665(.a(n2727), .O(n2730));
  inv1   g2666(.a(n2728), .O(n2731));
  nor2   g2667(.a(n2731), .b(n2730), .O(n2732));
  nor2   g2668(.a(n2732), .b(n2729), .O(n2733));
  inv1   g2669(.a(n2733), .O(n2734));
  nor2   g2670(.a(n2734), .b(n2726), .O(n2735));
  inv1   g2671(.a(n2726), .O(n2736));
  nor2   g2672(.a(n2733), .b(n2736), .O(n2737));
  nor2   g2673(.a(n2737), .b(n2735), .O(n2738));
  inv1   g2674(.a(n2738), .O(n2739));
  nor2   g2675(.a(n2739), .b(n2725), .O(n2740));
  inv1   g2676(.a(n2725), .O(n2741));
  nor2   g2677(.a(n2738), .b(n2741), .O(n2742));
  nor2   g2678(.a(n2742), .b(n2740), .O(n2743));
  inv1   g2679(.a(n2743), .O(n2744));
  nor2   g2680(.a(n2744), .b(n2724), .O(n2745));
  inv1   g2681(.a(n2724), .O(n2746));
  nor2   g2682(.a(n2743), .b(n2746), .O(n2747));
  nor2   g2683(.a(n2747), .b(n2745), .O(n2748));
  inv1   g2684(.a(n2748), .O(n2749));
  nor2   g2685(.a(n2749), .b(n2723), .O(n2750));
  inv1   g2686(.a(n2723), .O(n2751));
  nor2   g2687(.a(n2748), .b(n2751), .O(n2752));
  nor2   g2688(.a(n2752), .b(n2750), .O(n2753));
  inv1   g2689(.a(n2753), .O(n2754));
  nor2   g2690(.a(n2754), .b(n2722), .O(n2755));
  inv1   g2691(.a(n2722), .O(n2756));
  nor2   g2692(.a(n2753), .b(n2756), .O(n2757));
  nor2   g2693(.a(n2757), .b(n2755), .O(n2758));
  inv1   g2694(.a(n2758), .O(n2759));
  nor2   g2695(.a(n2759), .b(n2721), .O(n2760));
  inv1   g2696(.a(n2721), .O(n2761));
  nor2   g2697(.a(n2758), .b(n2761), .O(n2762));
  nor2   g2698(.a(n2762), .b(n2760), .O(n2763));
  inv1   g2699(.a(n2763), .O(n2764));
  nor2   g2700(.a(n2764), .b(n2720), .O(n2765));
  inv1   g2701(.a(n2720), .O(n2766));
  nor2   g2702(.a(n2763), .b(n2766), .O(n2767));
  nor2   g2703(.a(n2767), .b(n2765), .O(n2768));
  inv1   g2704(.a(n2768), .O(n2769));
  nor2   g2705(.a(n2769), .b(n2719), .O(n2770));
  inv1   g2706(.a(n2719), .O(n2771));
  nor2   g2707(.a(n2768), .b(n2771), .O(n2772));
  nor2   g2708(.a(n2772), .b(n2770), .O(n2773));
  inv1   g2709(.a(n2773), .O(n2774));
  nor2   g2710(.a(n2774), .b(n2718), .O(n2775));
  inv1   g2711(.a(n2718), .O(n2776));
  nor2   g2712(.a(n2773), .b(n2776), .O(n2777));
  nor2   g2713(.a(n2777), .b(n2775), .O(n2778));
  inv1   g2714(.a(n2778), .O(G6250gat));
  nor2   g2715(.a(n2775), .b(n2770), .O(n2780));
  nor2   g2716(.a(n2765), .b(n2760), .O(n2781));
  nor2   g2717(.a(n1275), .b(n842), .O(n2782));
  nor2   g2718(.a(n2755), .b(n2750), .O(n2783));
  nor2   g2719(.a(n1111), .b(n984), .O(n2784));
  nor2   g2720(.a(n2745), .b(n2740), .O(n2785));
  nor2   g2721(.a(n959), .b(n1138), .O(n2786));
  nor2   g2722(.a(n819), .b(n1304), .O(n2787));
  nor2   g2723(.a(n2735), .b(n2729), .O(n2788));
  nor2   g2724(.a(n2788), .b(n2787), .O(n2789));
  inv1   g2725(.a(n2787), .O(n2790));
  inv1   g2726(.a(n2788), .O(n2791));
  nor2   g2727(.a(n2791), .b(n2790), .O(n2792));
  nor2   g2728(.a(n2792), .b(n2789), .O(n2793));
  inv1   g2729(.a(n2793), .O(n2794));
  nor2   g2730(.a(n2794), .b(n2786), .O(n2795));
  inv1   g2731(.a(n2786), .O(n2796));
  nor2   g2732(.a(n2793), .b(n2796), .O(n2797));
  nor2   g2733(.a(n2797), .b(n2795), .O(n2798));
  inv1   g2734(.a(n2798), .O(n2799));
  nor2   g2735(.a(n2799), .b(n2785), .O(n2800));
  inv1   g2736(.a(n2785), .O(n2801));
  nor2   g2737(.a(n2798), .b(n2801), .O(n2802));
  nor2   g2738(.a(n2802), .b(n2800), .O(n2803));
  inv1   g2739(.a(n2803), .O(n2804));
  nor2   g2740(.a(n2804), .b(n2784), .O(n2805));
  inv1   g2741(.a(n2784), .O(n2806));
  nor2   g2742(.a(n2803), .b(n2806), .O(n2807));
  nor2   g2743(.a(n2807), .b(n2805), .O(n2808));
  inv1   g2744(.a(n2808), .O(n2809));
  nor2   g2745(.a(n2809), .b(n2783), .O(n2810));
  inv1   g2746(.a(n2783), .O(n2811));
  nor2   g2747(.a(n2808), .b(n2811), .O(n2812));
  nor2   g2748(.a(n2812), .b(n2810), .O(n2813));
  inv1   g2749(.a(n2813), .O(n2814));
  nor2   g2750(.a(n2814), .b(n2782), .O(n2815));
  inv1   g2751(.a(n2782), .O(n2816));
  nor2   g2752(.a(n2813), .b(n2816), .O(n2817));
  nor2   g2753(.a(n2817), .b(n2815), .O(n2818));
  inv1   g2754(.a(n2818), .O(n2819));
  nor2   g2755(.a(n2819), .b(n2781), .O(n2820));
  inv1   g2756(.a(n2781), .O(n2821));
  nor2   g2757(.a(n2818), .b(n2821), .O(n2822));
  nor2   g2758(.a(n2822), .b(n2820), .O(n2823));
  inv1   g2759(.a(n2823), .O(n2824));
  nor2   g2760(.a(n2824), .b(n2780), .O(n2825));
  inv1   g2761(.a(n2780), .O(n2826));
  nor2   g2762(.a(n2823), .b(n2826), .O(n2827));
  nor2   g2763(.a(n2827), .b(n2825), .O(n2828));
  inv1   g2764(.a(n2828), .O(G6260gat));
  nor2   g2765(.a(n2825), .b(n2820), .O(n2830));
  nor2   g2766(.a(n2815), .b(n2810), .O(n2831));
  nor2   g2767(.a(n1275), .b(n984), .O(n2832));
  nor2   g2768(.a(n2805), .b(n2800), .O(n2833));
  nor2   g2769(.a(n1111), .b(n1138), .O(n2834));
  nor2   g2770(.a(n959), .b(n1304), .O(n2835));
  nor2   g2771(.a(n2795), .b(n2789), .O(n2836));
  nor2   g2772(.a(n2836), .b(n2835), .O(n2837));
  inv1   g2773(.a(n2835), .O(n2838));
  inv1   g2774(.a(n2836), .O(n2839));
  nor2   g2775(.a(n2839), .b(n2838), .O(n2840));
  nor2   g2776(.a(n2840), .b(n2837), .O(n2841));
  inv1   g2777(.a(n2841), .O(n2842));
  nor2   g2778(.a(n2842), .b(n2834), .O(n2843));
  inv1   g2779(.a(n2834), .O(n2844));
  nor2   g2780(.a(n2841), .b(n2844), .O(n2845));
  nor2   g2781(.a(n2845), .b(n2843), .O(n2846));
  inv1   g2782(.a(n2846), .O(n2847));
  nor2   g2783(.a(n2847), .b(n2833), .O(n2848));
  inv1   g2784(.a(n2833), .O(n2849));
  nor2   g2785(.a(n2846), .b(n2849), .O(n2850));
  nor2   g2786(.a(n2850), .b(n2848), .O(n2851));
  inv1   g2787(.a(n2851), .O(n2852));
  nor2   g2788(.a(n2852), .b(n2832), .O(n2853));
  inv1   g2789(.a(n2832), .O(n2854));
  nor2   g2790(.a(n2851), .b(n2854), .O(n2855));
  nor2   g2791(.a(n2855), .b(n2853), .O(n2856));
  inv1   g2792(.a(n2856), .O(n2857));
  nor2   g2793(.a(n2857), .b(n2831), .O(n2858));
  inv1   g2794(.a(n2831), .O(n2859));
  nor2   g2795(.a(n2856), .b(n2859), .O(n2860));
  nor2   g2796(.a(n2860), .b(n2858), .O(n2861));
  inv1   g2797(.a(n2861), .O(n2862));
  nor2   g2798(.a(n2862), .b(n2830), .O(n2863));
  inv1   g2799(.a(n2830), .O(n2864));
  nor2   g2800(.a(n2861), .b(n2864), .O(n2865));
  nor2   g2801(.a(n2865), .b(n2863), .O(n2866));
  inv1   g2802(.a(n2866), .O(G6270gat));
  nor2   g2803(.a(n2863), .b(n2858), .O(n2868));
  nor2   g2804(.a(n2853), .b(n2848), .O(n2869));
  nor2   g2805(.a(n1275), .b(n1138), .O(n2870));
  nor2   g2806(.a(n1111), .b(n1304), .O(n2871));
  nor2   g2807(.a(n2843), .b(n2837), .O(n2872));
  nor2   g2808(.a(n2872), .b(n2871), .O(n2873));
  inv1   g2809(.a(n2871), .O(n2874));
  inv1   g2810(.a(n2872), .O(n2875));
  nor2   g2811(.a(n2875), .b(n2874), .O(n2876));
  nor2   g2812(.a(n2876), .b(n2873), .O(n2877));
  inv1   g2813(.a(n2877), .O(n2878));
  nor2   g2814(.a(n2878), .b(n2870), .O(n2879));
  inv1   g2815(.a(n2870), .O(n2880));
  nor2   g2816(.a(n2877), .b(n2880), .O(n2881));
  nor2   g2817(.a(n2881), .b(n2879), .O(n2882));
  inv1   g2818(.a(n2882), .O(n2883));
  nor2   g2819(.a(n2883), .b(n2869), .O(n2884));
  inv1   g2820(.a(n2869), .O(n2885));
  nor2   g2821(.a(n2882), .b(n2885), .O(n2886));
  nor2   g2822(.a(n2886), .b(n2884), .O(n2887));
  inv1   g2823(.a(n2887), .O(n2888));
  nor2   g2824(.a(n2888), .b(n2868), .O(n2889));
  inv1   g2825(.a(n2868), .O(n2890));
  nor2   g2826(.a(n2887), .b(n2890), .O(n2891));
  nor2   g2827(.a(n2891), .b(n2889), .O(n2892));
  inv1   g2828(.a(n2892), .O(G6280gat));
  nor2   g2829(.a(n1275), .b(n1304), .O(n2894));
  nor2   g2830(.a(n2879), .b(n2873), .O(n2895));
  nor2   g2831(.a(n2895), .b(n2894), .O(n2896));
  nor2   g2832(.a(n2889), .b(n2884), .O(n2897));
  inv1   g2833(.a(n2894), .O(n2898));
  inv1   g2834(.a(n2895), .O(n2899));
  nor2   g2835(.a(n2899), .b(n2898), .O(n2900));
  nor2   g2836(.a(n2900), .b(n2896), .O(n2901));
  inv1   g2837(.a(n2901), .O(n2902));
  nor2   g2838(.a(n2902), .b(n2897), .O(n2903));
  nor2   g2839(.a(n2903), .b(n2896), .O(G6287gat));
  inv1   g2840(.a(n2897), .O(n2905));
  nor2   g2841(.a(n2901), .b(n2905), .O(n2906));
  nor2   g2842(.a(n2906), .b(n2903), .O(n2907));
  inv1   g2843(.a(n2907), .O(G6288gat));
endmodule


