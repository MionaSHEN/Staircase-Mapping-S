// Benchmark "c1355_blif" written by ABC on Sun Mar 24 18:39:13 2019

module c1355_blif  ( 
    G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat,
    G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat,
    G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat,
    G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat,
    G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat,
    G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat,
    G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat,
    G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat,
    G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat,
    G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n443, n444, n445, n446, n447, n449, n450, n451,
    n452, n453, n455, n456, n457, n458, n459, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472, n474, n475, n476, n477, n478,
    n480, n481, n482, n483, n484, n486, n487, n488, n489, n490, n492, n493,
    n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n506,
    n507, n508, n509, n510, n512, n513, n514, n515, n516, n518, n519, n520,
    n521, n522, n524, n525, n526, n527, n528, n529, n530, n531, n532, n534,
    n535, n536, n537, n538, n540, n541, n542, n543, n544, n546, n547, n548,
    n549, n550, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n573, n574,
    n575, n576, n577, n579, n580, n581, n582, n583, n585, n586, n587, n588,
    n589, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n602,
    n603, n604, n605, n606, n608, n609, n610, n611, n612, n614, n615, n616,
    n617, n618, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n631, n632, n633, n634, n635, n637, n638, n639, n640, n641, n643, n644,
    n645, n646, n647, n649, n650, n651, n652, n653, n654, n655, n656, n657,
    n659, n660, n661, n662, n663, n665, n666, n667, n668, n669, n671, n672,
    n673, n674, n675;
  inv1   g000(.a(G1gat), .O(n74));
  inv1   g001(.a(G225gat), .O(n75));
  inv1   g002(.a(G233gat), .O(n76));
  nor2   g003(.a(n76), .b(n75), .O(n77));
  inv1   g004(.a(n77), .O(n78));
  nor2   g005(.a(G57gat), .b(G29gat), .O(n79));
  inv1   g006(.a(G29gat), .O(n80));
  inv1   g007(.a(G57gat), .O(n81));
  nor2   g008(.a(n81), .b(n80), .O(n82));
  nor2   g009(.a(n82), .b(n79), .O(n83));
  nor2   g010(.a(n83), .b(n78), .O(n84));
  inv1   g011(.a(n83), .O(n85));
  nor2   g012(.a(n85), .b(n77), .O(n86));
  nor2   g013(.a(n86), .b(n84), .O(n87));
  inv1   g014(.a(n87), .O(n88));
  nor2   g015(.a(G127gat), .b(G120gat), .O(n89));
  inv1   g016(.a(G120gat), .O(n90));
  inv1   g017(.a(G127gat), .O(n91));
  nor2   g018(.a(n91), .b(n90), .O(n92));
  nor2   g019(.a(n92), .b(n89), .O(n93));
  inv1   g020(.a(n93), .O(n94));
  inv1   g021(.a(G113gat), .O(n95));
  nor2   g022(.a(G134gat), .b(n95), .O(n96));
  inv1   g023(.a(G134gat), .O(n97));
  nor2   g024(.a(n97), .b(G113gat), .O(n98));
  nor2   g025(.a(n98), .b(n96), .O(n99));
  inv1   g026(.a(n99), .O(n100));
  nor2   g027(.a(n100), .b(n94), .O(n101));
  nor2   g028(.a(n99), .b(n93), .O(n102));
  nor2   g029(.a(n102), .b(n101), .O(n103));
  nor2   g030(.a(G155gat), .b(G148gat), .O(n104));
  inv1   g031(.a(G148gat), .O(n105));
  inv1   g032(.a(G155gat), .O(n106));
  nor2   g033(.a(n106), .b(n105), .O(n107));
  nor2   g034(.a(n107), .b(n104), .O(n108));
  inv1   g035(.a(n108), .O(n109));
  inv1   g036(.a(G141gat), .O(n110));
  nor2   g037(.a(G162gat), .b(n110), .O(n111));
  inv1   g038(.a(G162gat), .O(n112));
  nor2   g039(.a(n112), .b(G141gat), .O(n113));
  nor2   g040(.a(n113), .b(n111), .O(n114));
  inv1   g041(.a(n114), .O(n115));
  nor2   g042(.a(n115), .b(n109), .O(n116));
  nor2   g043(.a(n114), .b(n108), .O(n117));
  nor2   g044(.a(n117), .b(n116), .O(n118));
  inv1   g045(.a(n118), .O(n119));
  nor2   g046(.a(G85gat), .b(n74), .O(n120));
  inv1   g047(.a(G85gat), .O(n121));
  nor2   g048(.a(n121), .b(G1gat), .O(n122));
  nor2   g049(.a(n122), .b(n120), .O(n123));
  inv1   g050(.a(n123), .O(n124));
  nor2   g051(.a(n124), .b(n119), .O(n125));
  nor2   g052(.a(n123), .b(n118), .O(n126));
  nor2   g053(.a(n126), .b(n125), .O(n127));
  inv1   g054(.a(n127), .O(n128));
  nor2   g055(.a(n128), .b(n103), .O(n129));
  inv1   g056(.a(n103), .O(n130));
  nor2   g057(.a(n127), .b(n130), .O(n131));
  nor2   g058(.a(n131), .b(n129), .O(n132));
  inv1   g059(.a(n132), .O(n133));
  nor2   g060(.a(n133), .b(n88), .O(n134));
  nor2   g061(.a(n132), .b(n87), .O(n135));
  nor2   g062(.a(n135), .b(n134), .O(n136));
  inv1   g063(.a(G50gat), .O(n137));
  inv1   g064(.a(G22gat), .O(n138));
  inv1   g065(.a(G197gat), .O(n139));
  nor2   g066(.a(G218gat), .b(n139), .O(n140));
  inv1   g067(.a(G218gat), .O(n141));
  nor2   g068(.a(n141), .b(G197gat), .O(n142));
  nor2   g069(.a(n142), .b(n140), .O(n143));
  inv1   g070(.a(n143), .O(n144));
  inv1   g071(.a(G204gat), .O(n145));
  nor2   g072(.a(G211gat), .b(n145), .O(n146));
  inv1   g073(.a(G211gat), .O(n147));
  nor2   g074(.a(n147), .b(G204gat), .O(n148));
  nor2   g075(.a(n148), .b(n146), .O(n149));
  inv1   g076(.a(n149), .O(n150));
  nor2   g077(.a(n150), .b(n144), .O(n151));
  nor2   g078(.a(n149), .b(n143), .O(n152));
  nor2   g079(.a(n152), .b(n151), .O(n153));
  nor2   g080(.a(n153), .b(n138), .O(n154));
  inv1   g081(.a(n153), .O(n155));
  nor2   g082(.a(n155), .b(G22gat), .O(n156));
  nor2   g083(.a(n156), .b(n154), .O(n157));
  inv1   g084(.a(n157), .O(n158));
  nor2   g085(.a(n158), .b(n137), .O(n159));
  nor2   g086(.a(n157), .b(G50gat), .O(n160));
  nor2   g087(.a(n160), .b(n159), .O(n161));
  inv1   g088(.a(n161), .O(n162));
  inv1   g089(.a(G78gat), .O(n163));
  nor2   g090(.a(G106gat), .b(n163), .O(n164));
  inv1   g091(.a(G106gat), .O(n165));
  nor2   g092(.a(n165), .b(G78gat), .O(n166));
  nor2   g093(.a(n166), .b(n164), .O(n167));
  inv1   g094(.a(n167), .O(n168));
  inv1   g095(.a(G228gat), .O(n169));
  nor2   g096(.a(n76), .b(n169), .O(n170));
  inv1   g097(.a(n170), .O(n171));
  nor2   g098(.a(n171), .b(n118), .O(n172));
  nor2   g099(.a(n170), .b(n119), .O(n173));
  nor2   g100(.a(n173), .b(n172), .O(n174));
  nor2   g101(.a(n174), .b(n168), .O(n175));
  inv1   g102(.a(n174), .O(n176));
  nor2   g103(.a(n176), .b(n167), .O(n177));
  nor2   g104(.a(n177), .b(n175), .O(n178));
  inv1   g105(.a(n178), .O(n179));
  nor2   g106(.a(n179), .b(n162), .O(n180));
  nor2   g107(.a(n178), .b(n161), .O(n181));
  nor2   g108(.a(n181), .b(n180), .O(n182));
  inv1   g109(.a(G43gat), .O(n183));
  inv1   g110(.a(G15gat), .O(n184));
  inv1   g111(.a(G169gat), .O(n185));
  nor2   g112(.a(G190gat), .b(n185), .O(n186));
  inv1   g113(.a(G190gat), .O(n187));
  nor2   g114(.a(n187), .b(G169gat), .O(n188));
  nor2   g115(.a(n188), .b(n186), .O(n189));
  inv1   g116(.a(n189), .O(n190));
  inv1   g117(.a(G176gat), .O(n191));
  nor2   g118(.a(G183gat), .b(n191), .O(n192));
  inv1   g119(.a(G183gat), .O(n193));
  nor2   g120(.a(n193), .b(G176gat), .O(n194));
  nor2   g121(.a(n194), .b(n192), .O(n195));
  inv1   g122(.a(n195), .O(n196));
  nor2   g123(.a(n196), .b(n190), .O(n197));
  nor2   g124(.a(n195), .b(n189), .O(n198));
  nor2   g125(.a(n198), .b(n197), .O(n199));
  nor2   g126(.a(n199), .b(n184), .O(n200));
  inv1   g127(.a(n199), .O(n201));
  nor2   g128(.a(n201), .b(G15gat), .O(n202));
  nor2   g129(.a(n202), .b(n200), .O(n203));
  inv1   g130(.a(n203), .O(n204));
  nor2   g131(.a(n204), .b(n183), .O(n205));
  nor2   g132(.a(n203), .b(G43gat), .O(n206));
  nor2   g133(.a(n206), .b(n205), .O(n207));
  inv1   g134(.a(n207), .O(n208));
  inv1   g135(.a(G71gat), .O(n209));
  nor2   g136(.a(G99gat), .b(n209), .O(n210));
  inv1   g137(.a(G99gat), .O(n211));
  nor2   g138(.a(n211), .b(G71gat), .O(n212));
  nor2   g139(.a(n212), .b(n210), .O(n213));
  inv1   g140(.a(n213), .O(n214));
  inv1   g141(.a(G227gat), .O(n215));
  nor2   g142(.a(n76), .b(n215), .O(n216));
  inv1   g143(.a(n216), .O(n217));
  nor2   g144(.a(n217), .b(n103), .O(n218));
  nor2   g145(.a(n216), .b(n130), .O(n219));
  nor2   g146(.a(n219), .b(n218), .O(n220));
  nor2   g147(.a(n220), .b(n214), .O(n221));
  inv1   g148(.a(n220), .O(n222));
  nor2   g149(.a(n222), .b(n213), .O(n223));
  nor2   g150(.a(n223), .b(n221), .O(n224));
  inv1   g151(.a(n224), .O(n225));
  nor2   g152(.a(n225), .b(n208), .O(n226));
  nor2   g153(.a(n224), .b(n207), .O(n227));
  nor2   g154(.a(n227), .b(n226), .O(n228));
  inv1   g155(.a(n228), .O(n229));
  nor2   g156(.a(n229), .b(n182), .O(n230));
  inv1   g157(.a(n182), .O(n231));
  nor2   g158(.a(n228), .b(n231), .O(n232));
  nor2   g159(.a(n232), .b(n230), .O(n233));
  inv1   g160(.a(n136), .O(n234));
  inv1   g161(.a(G64gat), .O(n235));
  nor2   g162(.a(G92gat), .b(n235), .O(n236));
  inv1   g163(.a(G92gat), .O(n237));
  nor2   g164(.a(n237), .b(G64gat), .O(n238));
  nor2   g165(.a(n238), .b(n236), .O(n239));
  inv1   g166(.a(n239), .O(n240));
  nor2   g167(.a(n240), .b(n199), .O(n241));
  nor2   g168(.a(n239), .b(n201), .O(n242));
  nor2   g169(.a(n242), .b(n241), .O(n243));
  inv1   g170(.a(n243), .O(n244));
  inv1   g171(.a(G226gat), .O(n245));
  nor2   g172(.a(n76), .b(n245), .O(n246));
  inv1   g173(.a(n246), .O(n247));
  nor2   g174(.a(n247), .b(n155), .O(n248));
  nor2   g175(.a(n246), .b(n153), .O(n249));
  nor2   g176(.a(n249), .b(n248), .O(n250));
  inv1   g177(.a(n250), .O(n251));
  inv1   g178(.a(G8gat), .O(n252));
  nor2   g179(.a(G36gat), .b(n252), .O(n253));
  inv1   g180(.a(G36gat), .O(n254));
  nor2   g181(.a(n254), .b(G8gat), .O(n255));
  nor2   g182(.a(n255), .b(n253), .O(n256));
  nor2   g183(.a(n256), .b(n251), .O(n257));
  inv1   g184(.a(n256), .O(n258));
  nor2   g185(.a(n258), .b(n250), .O(n259));
  nor2   g186(.a(n259), .b(n257), .O(n260));
  inv1   g187(.a(n260), .O(n261));
  nor2   g188(.a(n261), .b(n244), .O(n262));
  nor2   g189(.a(n260), .b(n243), .O(n263));
  nor2   g190(.a(n263), .b(n262), .O(n264));
  nor2   g191(.a(n264), .b(n234), .O(n265));
  inv1   g192(.a(n265), .O(n266));
  nor2   g193(.a(n266), .b(n233), .O(n267));
  inv1   g194(.a(n264), .O(n268));
  nor2   g195(.a(n268), .b(n234), .O(n269));
  nor2   g196(.a(n264), .b(n136), .O(n270));
  nor2   g197(.a(n270), .b(n269), .O(n271));
  nor2   g198(.a(n229), .b(n231), .O(n272));
  inv1   g199(.a(n272), .O(n273));
  nor2   g200(.a(n273), .b(n271), .O(n274));
  nor2   g201(.a(n274), .b(n267), .O(n275));
  inv1   g202(.a(G229gat), .O(n276));
  nor2   g203(.a(n76), .b(n276), .O(n277));
  inv1   g204(.a(n277), .O(n278));
  nor2   g205(.a(G141gat), .b(G113gat), .O(n279));
  nor2   g206(.a(n110), .b(n95), .O(n280));
  nor2   g207(.a(n280), .b(n279), .O(n281));
  nor2   g208(.a(n281), .b(n278), .O(n282));
  inv1   g209(.a(n281), .O(n283));
  nor2   g210(.a(n283), .b(n277), .O(n284));
  nor2   g211(.a(n284), .b(n282), .O(n285));
  inv1   g212(.a(n285), .O(n286));
  nor2   g213(.a(G197gat), .b(n185), .O(n287));
  nor2   g214(.a(n139), .b(G169gat), .O(n288));
  nor2   g215(.a(n288), .b(n287), .O(n289));
  inv1   g216(.a(n289), .O(n290));
  nor2   g217(.a(G15gat), .b(G8gat), .O(n291));
  nor2   g218(.a(n184), .b(n252), .O(n292));
  nor2   g219(.a(n292), .b(n291), .O(n293));
  inv1   g220(.a(n293), .O(n294));
  nor2   g221(.a(G22gat), .b(n74), .O(n295));
  nor2   g222(.a(n138), .b(G1gat), .O(n296));
  nor2   g223(.a(n296), .b(n295), .O(n297));
  inv1   g224(.a(n297), .O(n298));
  nor2   g225(.a(n298), .b(n294), .O(n299));
  nor2   g226(.a(n297), .b(n293), .O(n300));
  nor2   g227(.a(n300), .b(n299), .O(n301));
  inv1   g228(.a(n301), .O(n302));
  nor2   g229(.a(n302), .b(n290), .O(n303));
  nor2   g230(.a(n301), .b(n289), .O(n304));
  nor2   g231(.a(n304), .b(n303), .O(n305));
  inv1   g232(.a(n305), .O(n306));
  nor2   g233(.a(G43gat), .b(G36gat), .O(n307));
  nor2   g234(.a(n183), .b(n254), .O(n308));
  nor2   g235(.a(n308), .b(n307), .O(n309));
  inv1   g236(.a(n309), .O(n310));
  nor2   g237(.a(G50gat), .b(n80), .O(n311));
  nor2   g238(.a(n137), .b(G29gat), .O(n312));
  nor2   g239(.a(n312), .b(n311), .O(n313));
  inv1   g240(.a(n313), .O(n314));
  nor2   g241(.a(n314), .b(n310), .O(n315));
  nor2   g242(.a(n313), .b(n309), .O(n316));
  nor2   g243(.a(n316), .b(n315), .O(n317));
  nor2   g244(.a(n317), .b(n306), .O(n318));
  inv1   g245(.a(n317), .O(n319));
  nor2   g246(.a(n319), .b(n305), .O(n320));
  nor2   g247(.a(n320), .b(n318), .O(n321));
  inv1   g248(.a(n321), .O(n322));
  nor2   g249(.a(n322), .b(n286), .O(n323));
  nor2   g250(.a(n321), .b(n285), .O(n324));
  nor2   g251(.a(n324), .b(n323), .O(n325));
  nor2   g252(.a(G204gat), .b(n191), .O(n326));
  nor2   g253(.a(n145), .b(G176gat), .O(n327));
  nor2   g254(.a(n327), .b(n326), .O(n328));
  inv1   g255(.a(n328), .O(n329));
  nor2   g256(.a(G78gat), .b(n81), .O(n330));
  nor2   g257(.a(n163), .b(G57gat), .O(n331));
  nor2   g258(.a(n331), .b(n330), .O(n332));
  inv1   g259(.a(n332), .O(n333));
  nor2   g260(.a(G71gat), .b(n235), .O(n334));
  nor2   g261(.a(n209), .b(G64gat), .O(n335));
  nor2   g262(.a(n335), .b(n334), .O(n336));
  inv1   g263(.a(n336), .O(n337));
  nor2   g264(.a(n337), .b(n333), .O(n338));
  nor2   g265(.a(n336), .b(n332), .O(n339));
  nor2   g266(.a(n339), .b(n338), .O(n340));
  nor2   g267(.a(n340), .b(n329), .O(n341));
  inv1   g268(.a(n340), .O(n342));
  nor2   g269(.a(n342), .b(n328), .O(n343));
  nor2   g270(.a(n343), .b(n341), .O(n344));
  inv1   g271(.a(n344), .O(n345));
  inv1   g272(.a(G230gat), .O(n346));
  nor2   g273(.a(n76), .b(n346), .O(n347));
  inv1   g274(.a(n347), .O(n348));
  nor2   g275(.a(G106gat), .b(n121), .O(n349));
  nor2   g276(.a(n165), .b(G85gat), .O(n350));
  nor2   g277(.a(n350), .b(n349), .O(n351));
  inv1   g278(.a(n351), .O(n352));
  nor2   g279(.a(G99gat), .b(n237), .O(n353));
  nor2   g280(.a(n211), .b(G92gat), .O(n354));
  nor2   g281(.a(n354), .b(n353), .O(n355));
  inv1   g282(.a(n355), .O(n356));
  nor2   g283(.a(n356), .b(n352), .O(n357));
  nor2   g284(.a(n355), .b(n351), .O(n358));
  nor2   g285(.a(n358), .b(n357), .O(n359));
  inv1   g286(.a(n359), .O(n360));
  nor2   g287(.a(n360), .b(n348), .O(n361));
  nor2   g288(.a(n359), .b(n347), .O(n362));
  nor2   g289(.a(n362), .b(n361), .O(n363));
  inv1   g290(.a(n363), .O(n364));
  nor2   g291(.a(G148gat), .b(n90), .O(n365));
  nor2   g292(.a(n105), .b(G120gat), .O(n366));
  nor2   g293(.a(n366), .b(n365), .O(n367));
  nor2   g294(.a(n367), .b(n364), .O(n368));
  inv1   g295(.a(n367), .O(n369));
  nor2   g296(.a(n369), .b(n363), .O(n370));
  nor2   g297(.a(n370), .b(n368), .O(n371));
  inv1   g298(.a(n371), .O(n372));
  nor2   g299(.a(n372), .b(n345), .O(n373));
  nor2   g300(.a(n371), .b(n344), .O(n374));
  nor2   g301(.a(n374), .b(n373), .O(n375));
  nor2   g302(.a(n375), .b(n325), .O(n376));
  inv1   g303(.a(n376), .O(n377));
  nor2   g304(.a(n359), .b(n97), .O(n378));
  nor2   g305(.a(n360), .b(G134gat), .O(n379));
  nor2   g306(.a(n379), .b(n378), .O(n380));
  inv1   g307(.a(n380), .O(n381));
  nor2   g308(.a(n381), .b(n112), .O(n382));
  nor2   g309(.a(n380), .b(G162gat), .O(n383));
  nor2   g310(.a(n383), .b(n382), .O(n384));
  inv1   g311(.a(n384), .O(n385));
  nor2   g312(.a(G218gat), .b(n187), .O(n386));
  nor2   g313(.a(n141), .b(G190gat), .O(n387));
  nor2   g314(.a(n387), .b(n386), .O(n388));
  inv1   g315(.a(n388), .O(n389));
  inv1   g316(.a(G232gat), .O(n390));
  nor2   g317(.a(n76), .b(n390), .O(n391));
  inv1   g318(.a(n391), .O(n392));
  nor2   g319(.a(n392), .b(n317), .O(n393));
  nor2   g320(.a(n391), .b(n319), .O(n394));
  nor2   g321(.a(n394), .b(n393), .O(n395));
  nor2   g322(.a(n395), .b(n389), .O(n396));
  inv1   g323(.a(n395), .O(n397));
  nor2   g324(.a(n397), .b(n388), .O(n398));
  nor2   g325(.a(n398), .b(n396), .O(n399));
  inv1   g326(.a(n399), .O(n400));
  nor2   g327(.a(n400), .b(n385), .O(n401));
  nor2   g328(.a(n399), .b(n384), .O(n402));
  nor2   g329(.a(n402), .b(n401), .O(n403));
  inv1   g330(.a(n403), .O(n404));
  nor2   g331(.a(n340), .b(n91), .O(n405));
  nor2   g332(.a(n342), .b(G127gat), .O(n406));
  nor2   g333(.a(n406), .b(n405), .O(n407));
  inv1   g334(.a(n407), .O(n408));
  nor2   g335(.a(n408), .b(n106), .O(n409));
  nor2   g336(.a(n407), .b(G155gat), .O(n410));
  nor2   g337(.a(n410), .b(n409), .O(n411));
  inv1   g338(.a(n411), .O(n412));
  nor2   g339(.a(G211gat), .b(n193), .O(n413));
  nor2   g340(.a(n147), .b(G183gat), .O(n414));
  nor2   g341(.a(n414), .b(n413), .O(n415));
  inv1   g342(.a(n415), .O(n416));
  inv1   g343(.a(G231gat), .O(n417));
  nor2   g344(.a(n76), .b(n417), .O(n418));
  inv1   g345(.a(n418), .O(n419));
  nor2   g346(.a(n419), .b(n301), .O(n420));
  nor2   g347(.a(n418), .b(n302), .O(n421));
  nor2   g348(.a(n421), .b(n420), .O(n422));
  nor2   g349(.a(n422), .b(n416), .O(n423));
  inv1   g350(.a(n422), .O(n424));
  nor2   g351(.a(n424), .b(n415), .O(n425));
  nor2   g352(.a(n425), .b(n423), .O(n426));
  inv1   g353(.a(n426), .O(n427));
  nor2   g354(.a(n427), .b(n412), .O(n428));
  nor2   g355(.a(n426), .b(n411), .O(n429));
  nor2   g356(.a(n429), .b(n428), .O(n430));
  nor2   g357(.a(n430), .b(n404), .O(n431));
  inv1   g358(.a(n431), .O(n432));
  nor2   g359(.a(n432), .b(n377), .O(n433));
  inv1   g360(.a(n433), .O(n434));
  nor2   g361(.a(n434), .b(n275), .O(n435));
  inv1   g362(.a(n435), .O(n436));
  nor2   g363(.a(n436), .b(n136), .O(n437));
  nor2   g364(.a(n437), .b(n74), .O(n438));
  inv1   g365(.a(n437), .O(n439));
  nor2   g366(.a(n439), .b(G1gat), .O(n440));
  nor2   g367(.a(n440), .b(n438), .O(n441));
  inv1   g368(.a(n441), .O(G1324gat));
  nor2   g369(.a(n436), .b(n268), .O(n443));
  nor2   g370(.a(n443), .b(n252), .O(n444));
  inv1   g371(.a(n443), .O(n445));
  nor2   g372(.a(n445), .b(G8gat), .O(n446));
  nor2   g373(.a(n446), .b(n444), .O(n447));
  inv1   g374(.a(n447), .O(G1325gat));
  nor2   g375(.a(n436), .b(n228), .O(n449));
  nor2   g376(.a(n449), .b(n184), .O(n450));
  inv1   g377(.a(n449), .O(n451));
  nor2   g378(.a(n451), .b(G15gat), .O(n452));
  nor2   g379(.a(n452), .b(n450), .O(n453));
  inv1   g380(.a(n453), .O(G1326gat));
  nor2   g381(.a(n436), .b(n182), .O(n455));
  nor2   g382(.a(n455), .b(n138), .O(n456));
  inv1   g383(.a(n455), .O(n457));
  nor2   g384(.a(n457), .b(G22gat), .O(n458));
  nor2   g385(.a(n458), .b(n456), .O(n459));
  inv1   g386(.a(n459), .O(G1327gat));
  inv1   g387(.a(n430), .O(n461));
  nor2   g388(.a(n461), .b(n403), .O(n462));
  inv1   g389(.a(n462), .O(n463));
  nor2   g390(.a(n463), .b(n377), .O(n464));
  inv1   g391(.a(n464), .O(n465));
  nor2   g392(.a(n465), .b(n275), .O(n466));
  inv1   g393(.a(n466), .O(n467));
  nor2   g394(.a(n467), .b(n136), .O(n468));
  nor2   g395(.a(n468), .b(n80), .O(n469));
  inv1   g396(.a(n468), .O(n470));
  nor2   g397(.a(n470), .b(G29gat), .O(n471));
  nor2   g398(.a(n471), .b(n469), .O(n472));
  inv1   g399(.a(n472), .O(G1328gat));
  nor2   g400(.a(n467), .b(n268), .O(n474));
  nor2   g401(.a(n474), .b(n254), .O(n475));
  inv1   g402(.a(n474), .O(n476));
  nor2   g403(.a(n476), .b(G36gat), .O(n477));
  nor2   g404(.a(n477), .b(n475), .O(n478));
  inv1   g405(.a(n478), .O(G1329gat));
  nor2   g406(.a(n467), .b(n228), .O(n480));
  nor2   g407(.a(n480), .b(n183), .O(n481));
  inv1   g408(.a(n480), .O(n482));
  nor2   g409(.a(n482), .b(G43gat), .O(n483));
  nor2   g410(.a(n483), .b(n481), .O(n484));
  inv1   g411(.a(n484), .O(G1330gat));
  nor2   g412(.a(n467), .b(n182), .O(n486));
  nor2   g413(.a(n486), .b(n137), .O(n487));
  inv1   g414(.a(n486), .O(n488));
  nor2   g415(.a(n488), .b(G50gat), .O(n489));
  nor2   g416(.a(n489), .b(n487), .O(n490));
  inv1   g417(.a(n490), .O(G1331gat));
  inv1   g418(.a(n325), .O(n492));
  inv1   g419(.a(n375), .O(n493));
  nor2   g420(.a(n493), .b(n492), .O(n494));
  inv1   g421(.a(n494), .O(n495));
  nor2   g422(.a(n495), .b(n432), .O(n496));
  inv1   g423(.a(n496), .O(n497));
  nor2   g424(.a(n497), .b(n275), .O(n498));
  inv1   g425(.a(n498), .O(n499));
  nor2   g426(.a(n499), .b(n136), .O(n500));
  nor2   g427(.a(n500), .b(n81), .O(n501));
  inv1   g428(.a(n500), .O(n502));
  nor2   g429(.a(n502), .b(G57gat), .O(n503));
  nor2   g430(.a(n503), .b(n501), .O(n504));
  inv1   g431(.a(n504), .O(G1332gat));
  nor2   g432(.a(n499), .b(n268), .O(n506));
  nor2   g433(.a(n506), .b(n235), .O(n507));
  inv1   g434(.a(n506), .O(n508));
  nor2   g435(.a(n508), .b(G64gat), .O(n509));
  nor2   g436(.a(n509), .b(n507), .O(n510));
  inv1   g437(.a(n510), .O(G1333gat));
  nor2   g438(.a(n499), .b(n228), .O(n512));
  nor2   g439(.a(n512), .b(n209), .O(n513));
  inv1   g440(.a(n512), .O(n514));
  nor2   g441(.a(n514), .b(G71gat), .O(n515));
  nor2   g442(.a(n515), .b(n513), .O(n516));
  inv1   g443(.a(n516), .O(G1334gat));
  nor2   g444(.a(n499), .b(n182), .O(n518));
  nor2   g445(.a(n518), .b(n163), .O(n519));
  inv1   g446(.a(n518), .O(n520));
  nor2   g447(.a(n520), .b(G78gat), .O(n521));
  nor2   g448(.a(n521), .b(n519), .O(n522));
  inv1   g449(.a(n522), .O(G1335gat));
  nor2   g450(.a(n495), .b(n463), .O(n524));
  inv1   g451(.a(n524), .O(n525));
  nor2   g452(.a(n525), .b(n275), .O(n526));
  inv1   g453(.a(n526), .O(n527));
  nor2   g454(.a(n527), .b(n136), .O(n528));
  nor2   g455(.a(n528), .b(n121), .O(n529));
  inv1   g456(.a(n528), .O(n530));
  nor2   g457(.a(n530), .b(G85gat), .O(n531));
  nor2   g458(.a(n531), .b(n529), .O(n532));
  inv1   g459(.a(n532), .O(G1336gat));
  nor2   g460(.a(n527), .b(n268), .O(n534));
  nor2   g461(.a(n534), .b(n237), .O(n535));
  inv1   g462(.a(n534), .O(n536));
  nor2   g463(.a(n536), .b(G92gat), .O(n537));
  nor2   g464(.a(n537), .b(n535), .O(n538));
  inv1   g465(.a(n538), .O(G1337gat));
  nor2   g466(.a(n527), .b(n228), .O(n540));
  nor2   g467(.a(n540), .b(n211), .O(n541));
  inv1   g468(.a(n540), .O(n542));
  nor2   g469(.a(n542), .b(G99gat), .O(n543));
  nor2   g470(.a(n543), .b(n541), .O(n544));
  inv1   g471(.a(n544), .O(G1338gat));
  nor2   g472(.a(n527), .b(n182), .O(n546));
  nor2   g473(.a(n546), .b(n165), .O(n547));
  inv1   g474(.a(n546), .O(n548));
  nor2   g475(.a(n548), .b(G106gat), .O(n549));
  nor2   g476(.a(n549), .b(n547), .O(n550));
  inv1   g477(.a(n550), .O(G1339gat));
  nor2   g478(.a(n462), .b(n431), .O(n552));
  nor2   g479(.a(n375), .b(n492), .O(n553));
  inv1   g480(.a(n553), .O(n554));
  nor2   g481(.a(n554), .b(n552), .O(n555));
  nor2   g482(.a(n494), .b(n376), .O(n556));
  nor2   g483(.a(n461), .b(n404), .O(n557));
  inv1   g484(.a(n557), .O(n558));
  nor2   g485(.a(n558), .b(n556), .O(n559));
  nor2   g486(.a(n559), .b(n555), .O(n560));
  inv1   g487(.a(n232), .O(n561));
  inv1   g488(.a(n270), .O(n562));
  nor2   g489(.a(n562), .b(n561), .O(n563));
  inv1   g490(.a(n563), .O(n564));
  nor2   g491(.a(n564), .b(n560), .O(n565));
  inv1   g492(.a(n565), .O(n566));
  nor2   g493(.a(n566), .b(n325), .O(n567));
  nor2   g494(.a(n567), .b(n95), .O(n568));
  inv1   g495(.a(n567), .O(n569));
  nor2   g496(.a(n569), .b(G113gat), .O(n570));
  nor2   g497(.a(n570), .b(n568), .O(n571));
  inv1   g498(.a(n571), .O(G1340gat));
  nor2   g499(.a(n566), .b(n493), .O(n573));
  nor2   g500(.a(n573), .b(n90), .O(n574));
  inv1   g501(.a(n573), .O(n575));
  nor2   g502(.a(n575), .b(G120gat), .O(n576));
  nor2   g503(.a(n576), .b(n574), .O(n577));
  inv1   g504(.a(n577), .O(G1341gat));
  nor2   g505(.a(n566), .b(n430), .O(n579));
  nor2   g506(.a(n579), .b(n91), .O(n580));
  inv1   g507(.a(n579), .O(n581));
  nor2   g508(.a(n581), .b(G127gat), .O(n582));
  nor2   g509(.a(n582), .b(n580), .O(n583));
  inv1   g510(.a(n583), .O(G1342gat));
  nor2   g511(.a(n566), .b(n403), .O(n585));
  nor2   g512(.a(n585), .b(n97), .O(n586));
  inv1   g513(.a(n585), .O(n587));
  nor2   g514(.a(n587), .b(G134gat), .O(n588));
  nor2   g515(.a(n588), .b(n586), .O(n589));
  inv1   g516(.a(n589), .O(G1343gat));
  inv1   g517(.a(n230), .O(n591));
  nor2   g518(.a(n562), .b(n591), .O(n592));
  inv1   g519(.a(n592), .O(n593));
  nor2   g520(.a(n593), .b(n560), .O(n594));
  inv1   g521(.a(n594), .O(n595));
  nor2   g522(.a(n595), .b(n325), .O(n596));
  nor2   g523(.a(n596), .b(n110), .O(n597));
  inv1   g524(.a(n596), .O(n598));
  nor2   g525(.a(n598), .b(G141gat), .O(n599));
  nor2   g526(.a(n599), .b(n597), .O(n600));
  inv1   g527(.a(n600), .O(G1344gat));
  nor2   g528(.a(n595), .b(n493), .O(n602));
  nor2   g529(.a(n602), .b(n105), .O(n603));
  inv1   g530(.a(n602), .O(n604));
  nor2   g531(.a(n604), .b(G148gat), .O(n605));
  nor2   g532(.a(n605), .b(n603), .O(n606));
  inv1   g533(.a(n606), .O(G1345gat));
  nor2   g534(.a(n595), .b(n430), .O(n608));
  nor2   g535(.a(n608), .b(n106), .O(n609));
  inv1   g536(.a(n608), .O(n610));
  nor2   g537(.a(n610), .b(G155gat), .O(n611));
  nor2   g538(.a(n611), .b(n609), .O(n612));
  inv1   g539(.a(n612), .O(G1346gat));
  nor2   g540(.a(n595), .b(n403), .O(n614));
  nor2   g541(.a(n614), .b(n112), .O(n615));
  inv1   g542(.a(n614), .O(n616));
  nor2   g543(.a(n616), .b(G162gat), .O(n617));
  nor2   g544(.a(n617), .b(n615), .O(n618));
  inv1   g545(.a(n618), .O(G1347gat));
  inv1   g546(.a(n269), .O(n620));
  nor2   g547(.a(n620), .b(n561), .O(n621));
  inv1   g548(.a(n621), .O(n622));
  nor2   g549(.a(n622), .b(n560), .O(n623));
  inv1   g550(.a(n623), .O(n624));
  nor2   g551(.a(n624), .b(n325), .O(n625));
  nor2   g552(.a(n625), .b(n185), .O(n626));
  inv1   g553(.a(n625), .O(n627));
  nor2   g554(.a(n627), .b(G169gat), .O(n628));
  nor2   g555(.a(n628), .b(n626), .O(n629));
  inv1   g556(.a(n629), .O(G1348gat));
  nor2   g557(.a(n624), .b(n493), .O(n631));
  nor2   g558(.a(n631), .b(n191), .O(n632));
  inv1   g559(.a(n631), .O(n633));
  nor2   g560(.a(n633), .b(G176gat), .O(n634));
  nor2   g561(.a(n634), .b(n632), .O(n635));
  inv1   g562(.a(n635), .O(G1349gat));
  nor2   g563(.a(n624), .b(n430), .O(n637));
  nor2   g564(.a(n637), .b(n193), .O(n638));
  inv1   g565(.a(n637), .O(n639));
  nor2   g566(.a(n639), .b(G183gat), .O(n640));
  nor2   g567(.a(n640), .b(n638), .O(n641));
  inv1   g568(.a(n641), .O(G1350gat));
  nor2   g569(.a(n624), .b(n403), .O(n643));
  nor2   g570(.a(n643), .b(n187), .O(n644));
  inv1   g571(.a(n643), .O(n645));
  nor2   g572(.a(n645), .b(G190gat), .O(n646));
  nor2   g573(.a(n646), .b(n644), .O(n647));
  inv1   g574(.a(n647), .O(G1351gat));
  nor2   g575(.a(n620), .b(n591), .O(n649));
  inv1   g576(.a(n649), .O(n650));
  nor2   g577(.a(n650), .b(n560), .O(n651));
  inv1   g578(.a(n651), .O(n652));
  nor2   g579(.a(n652), .b(n325), .O(n653));
  nor2   g580(.a(n653), .b(n139), .O(n654));
  inv1   g581(.a(n653), .O(n655));
  nor2   g582(.a(n655), .b(G197gat), .O(n656));
  nor2   g583(.a(n656), .b(n654), .O(n657));
  inv1   g584(.a(n657), .O(G1352gat));
  nor2   g585(.a(n652), .b(n493), .O(n659));
  nor2   g586(.a(n659), .b(n145), .O(n660));
  inv1   g587(.a(n659), .O(n661));
  nor2   g588(.a(n661), .b(G204gat), .O(n662));
  nor2   g589(.a(n662), .b(n660), .O(n663));
  inv1   g590(.a(n663), .O(G1353gat));
  nor2   g591(.a(n652), .b(n430), .O(n665));
  nor2   g592(.a(n665), .b(n147), .O(n666));
  inv1   g593(.a(n665), .O(n667));
  nor2   g594(.a(n667), .b(G211gat), .O(n668));
  nor2   g595(.a(n668), .b(n666), .O(n669));
  inv1   g596(.a(n669), .O(G1354gat));
  nor2   g597(.a(n652), .b(n403), .O(n671));
  nor2   g598(.a(n671), .b(n141), .O(n672));
  inv1   g599(.a(n671), .O(n673));
  nor2   g600(.a(n673), .b(G218gat), .O(n674));
  nor2   g601(.a(n674), .b(n672), .O(n675));
  inv1   g602(.a(n675), .O(G1355gat));
endmodule


