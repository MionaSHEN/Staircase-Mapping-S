// Benchmark "c3540_blif" written by ABC on Sun Mar 24 18:39:14 2019

module c3540_blif  ( 
    G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
    G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200,
    G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274,
    G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698,
    G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107,
    G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
    G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270,
    G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire n73, n74, n75, n76, n78, n79, n80, n82, n83, n84, n85, n86, n87, n88,
    n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
    n163, n164, n165, n166, n167, n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592, n594, n595, n596, n597, n598,
    n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
    n611, n612, n613, n614, n615, n616, n617, n618, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
    n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
    n854, n855, n856, n857, n858, n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
    n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
    n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
    n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
    n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
    n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
    n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
    n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
    n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
    n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
    n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
    n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
    n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
    n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
    n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
    n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
    n1406, n1407, n1408, n1409, n1410, n1411, n1413, n1414, n1415, n1416,
    n1417, n1418, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
    n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1448,
    n1449, n1450;
  nor2   g0000(.a(G68), .b(G58), .O(n73));
  inv1   g0001(.a(n73), .O(n74));
  nor2   g0002(.a(n74), .b(G50), .O(n75));
  inv1   g0003(.a(n75), .O(n76));
  nor2   g0004(.a(n76), .b(G77), .O(G353));
  inv1   g0005(.a(G87), .O(n78));
  nor2   g0006(.a(G107), .b(G97), .O(n79));
  nor2   g0007(.a(n79), .b(n78), .O(n80));
  inv1   g0008(.a(n80), .O(G355));
  inv1   g0009(.a(G1), .O(n82));
  inv1   g0010(.a(G20), .O(n83));
  nor2   g0011(.a(n83), .b(n82), .O(n84));
  inv1   g0012(.a(G68), .O(n85));
  inv1   g0013(.a(G238), .O(n86));
  nor2   g0014(.a(n86), .b(n85), .O(n87));
  inv1   g0015(.a(G97), .O(n88));
  inv1   g0016(.a(G257), .O(n89));
  nor2   g0017(.a(n89), .b(n88), .O(n90));
  nor2   g0018(.a(n90), .b(n87), .O(n91));
  inv1   g0019(.a(n91), .O(n92));
  inv1   g0020(.a(G77), .O(n93));
  inv1   g0021(.a(G244), .O(n94));
  nor2   g0022(.a(n94), .b(n93), .O(n95));
  inv1   g0023(.a(G116), .O(n96));
  inv1   g0024(.a(G270), .O(n97));
  nor2   g0025(.a(n97), .b(n96), .O(n98));
  nor2   g0026(.a(n98), .b(n95), .O(n99));
  inv1   g0027(.a(n99), .O(n100));
  nor2   g0028(.a(n100), .b(n92), .O(n101));
  inv1   g0029(.a(n101), .O(n102));
  inv1   g0030(.a(G250), .O(n103));
  nor2   g0031(.a(n103), .b(n78), .O(n104));
  inv1   g0032(.a(G50), .O(n105));
  inv1   g0033(.a(G226), .O(n106));
  nor2   g0034(.a(n106), .b(n105), .O(n107));
  nor2   g0035(.a(n107), .b(n104), .O(n108));
  inv1   g0036(.a(n108), .O(n109));
  inv1   g0037(.a(G58), .O(n110));
  inv1   g0038(.a(G232), .O(n111));
  nor2   g0039(.a(n111), .b(n110), .O(n112));
  inv1   g0040(.a(G107), .O(n113));
  inv1   g0041(.a(G264), .O(n114));
  nor2   g0042(.a(n114), .b(n113), .O(n115));
  nor2   g0043(.a(n115), .b(n112), .O(n116));
  inv1   g0044(.a(n116), .O(n117));
  nor2   g0045(.a(n117), .b(n109), .O(n118));
  inv1   g0046(.a(n118), .O(n119));
  nor2   g0047(.a(n119), .b(n102), .O(n120));
  nor2   g0048(.a(n120), .b(n84), .O(n121));
  inv1   g0049(.a(G13), .O(n122));
  nor2   g0050(.a(n122), .b(n82), .O(n123));
  inv1   g0051(.a(n123), .O(n124));
  nor2   g0052(.a(n124), .b(n83), .O(n125));
  inv1   g0053(.a(n125), .O(n126));
  nor2   g0054(.a(n73), .b(n105), .O(n127));
  inv1   g0055(.a(n127), .O(n128));
  nor2   g0056(.a(n128), .b(n126), .O(n129));
  nor2   g0057(.a(G13), .b(n82), .O(n130));
  inv1   g0058(.a(n130), .O(n131));
  nor2   g0059(.a(n131), .b(n83), .O(n132));
  inv1   g0060(.a(n132), .O(n133));
  nor2   g0061(.a(G264), .b(G257), .O(n134));
  nor2   g0062(.a(n134), .b(n103), .O(n135));
  inv1   g0063(.a(n135), .O(n136));
  nor2   g0064(.a(n136), .b(n133), .O(n137));
  nor2   g0065(.a(n137), .b(n129), .O(n138));
  inv1   g0066(.a(n138), .O(n139));
  nor2   g0067(.a(n139), .b(n121), .O(G361));
  nor2   g0068(.a(G270), .b(n114), .O(n141));
  nor2   g0069(.a(n97), .b(G264), .O(n142));
  nor2   g0070(.a(n142), .b(n141), .O(n143));
  inv1   g0071(.a(n143), .O(n144));
  nor2   g0072(.a(G257), .b(n103), .O(n145));
  nor2   g0073(.a(n89), .b(G250), .O(n146));
  nor2   g0074(.a(n146), .b(n145), .O(n147));
  inv1   g0075(.a(n147), .O(n148));
  nor2   g0076(.a(n148), .b(n144), .O(n149));
  nor2   g0077(.a(n147), .b(n143), .O(n150));
  nor2   g0078(.a(n150), .b(n149), .O(n151));
  inv1   g0079(.a(n151), .O(n152));
  nor2   g0080(.a(G244), .b(n86), .O(n153));
  nor2   g0081(.a(n94), .b(G238), .O(n154));
  nor2   g0082(.a(n154), .b(n153), .O(n155));
  inv1   g0083(.a(n155), .O(n156));
  nor2   g0084(.a(G232), .b(n106), .O(n157));
  nor2   g0085(.a(n111), .b(G226), .O(n158));
  nor2   g0086(.a(n158), .b(n157), .O(n159));
  inv1   g0087(.a(n159), .O(n160));
  nor2   g0088(.a(n160), .b(n156), .O(n161));
  nor2   g0089(.a(n159), .b(n155), .O(n162));
  nor2   g0090(.a(n162), .b(n161), .O(n163));
  inv1   g0091(.a(n163), .O(n164));
  nor2   g0092(.a(n164), .b(n152), .O(n165));
  nor2   g0093(.a(n163), .b(n151), .O(n166));
  nor2   g0094(.a(n166), .b(n165), .O(n167));
  inv1   g0095(.a(n167), .O(G358));
  nor2   g0096(.a(n85), .b(n110), .O(n169));
  nor2   g0097(.a(n169), .b(n73), .O(n170));
  inv1   g0098(.a(n170), .O(n171));
  nor2   g0099(.a(n171), .b(n93), .O(n172));
  nor2   g0100(.a(n170), .b(G77), .O(n173));
  nor2   g0101(.a(n173), .b(n172), .O(n174));
  inv1   g0102(.a(n174), .O(n175));
  nor2   g0103(.a(n175), .b(n105), .O(n176));
  nor2   g0104(.a(n174), .b(G50), .O(n177));
  nor2   g0105(.a(n177), .b(n176), .O(n178));
  inv1   g0106(.a(n178), .O(n179));
  nor2   g0107(.a(n113), .b(n88), .O(n180));
  nor2   g0108(.a(n180), .b(n79), .O(n181));
  inv1   g0109(.a(n181), .O(n182));
  nor2   g0110(.a(G116), .b(n78), .O(n183));
  nor2   g0111(.a(n96), .b(G87), .O(n184));
  nor2   g0112(.a(n184), .b(n183), .O(n185));
  inv1   g0113(.a(n185), .O(n186));
  nor2   g0114(.a(n186), .b(n182), .O(n187));
  nor2   g0115(.a(n185), .b(n181), .O(n188));
  nor2   g0116(.a(n188), .b(n187), .O(n189));
  inv1   g0117(.a(n189), .O(n190));
  nor2   g0118(.a(n190), .b(n179), .O(n191));
  nor2   g0119(.a(n189), .b(n178), .O(n192));
  nor2   g0120(.a(n192), .b(n191), .O(G351));
  inv1   g0121(.a(G33), .O(n194));
  inv1   g0122(.a(G41), .O(n195));
  nor2   g0123(.a(n195), .b(n194), .O(n196));
  nor2   g0124(.a(n196), .b(n124), .O(n197));
  inv1   g0125(.a(n197), .O(n198));
  inv1   g0126(.a(G1698), .O(n199));
  nor2   g0127(.a(n199), .b(G33), .O(n200));
  inv1   g0128(.a(n200), .O(n201));
  nor2   g0129(.a(n201), .b(n94), .O(n202));
  nor2   g0130(.a(n96), .b(n194), .O(n203));
  nor2   g0131(.a(G1698), .b(G33), .O(n204));
  inv1   g0132(.a(n204), .O(n205));
  nor2   g0133(.a(n205), .b(n86), .O(n206));
  nor2   g0134(.a(n206), .b(n203), .O(n207));
  inv1   g0135(.a(n207), .O(n208));
  nor2   g0136(.a(n208), .b(n202), .O(n209));
  nor2   g0137(.a(n209), .b(n198), .O(n210));
  inv1   g0138(.a(G45), .O(n211));
  nor2   g0139(.a(n211), .b(G1), .O(n212));
  inv1   g0140(.a(n212), .O(n213));
  nor2   g0141(.a(n213), .b(G274), .O(n214));
  nor2   g0142(.a(n212), .b(G250), .O(n215));
  nor2   g0143(.a(n215), .b(n197), .O(n216));
  inv1   g0144(.a(n216), .O(n217));
  nor2   g0145(.a(n217), .b(n214), .O(n218));
  nor2   g0146(.a(n218), .b(n210), .O(n219));
  nor2   g0147(.a(n219), .b(G169), .O(n220));
  nor2   g0148(.a(n194), .b(G1), .O(n221));
  nor2   g0149(.a(n122), .b(G1), .O(n222));
  inv1   g0150(.a(n222), .O(n223));
  nor2   g0151(.a(n223), .b(n83), .O(n224));
  inv1   g0152(.a(n84), .O(n225));
  nor2   g0153(.a(n225), .b(n194), .O(n226));
  nor2   g0154(.a(n226), .b(n123), .O(n227));
  inv1   g0155(.a(n227), .O(n228));
  nor2   g0156(.a(n228), .b(n224), .O(n229));
  inv1   g0157(.a(n229), .O(n230));
  nor2   g0158(.a(n230), .b(n221), .O(n231));
  inv1   g0159(.a(n231), .O(n232));
  nor2   g0160(.a(n232), .b(n78), .O(n233));
  inv1   g0161(.a(n224), .O(n234));
  nor2   g0162(.a(n234), .b(G87), .O(n235));
  nor2   g0163(.a(n85), .b(G33), .O(n236));
  nor2   g0164(.a(n88), .b(n194), .O(n237));
  nor2   g0165(.a(n237), .b(G20), .O(n238));
  inv1   g0166(.a(n238), .O(n239));
  nor2   g0167(.a(n239), .b(n236), .O(n240));
  inv1   g0168(.a(n79), .O(n241));
  nor2   g0169(.a(n241), .b(G87), .O(n242));
  inv1   g0170(.a(n242), .O(n243));
  nor2   g0171(.a(n243), .b(n83), .O(n244));
  nor2   g0172(.a(n244), .b(n227), .O(n245));
  inv1   g0173(.a(n245), .O(n246));
  nor2   g0174(.a(n246), .b(n240), .O(n247));
  nor2   g0175(.a(n247), .b(n235), .O(n248));
  inv1   g0176(.a(n248), .O(n249));
  nor2   g0177(.a(n249), .b(n233), .O(n250));
  inv1   g0178(.a(n219), .O(n251));
  nor2   g0179(.a(n251), .b(G179), .O(n252));
  nor2   g0180(.a(n252), .b(n250), .O(n253));
  inv1   g0181(.a(n253), .O(n254));
  nor2   g0182(.a(n254), .b(n220), .O(n255));
  inv1   g0183(.a(n250), .O(n256));
  nor2   g0184(.a(n251), .b(G190), .O(n257));
  nor2   g0185(.a(n219), .b(G200), .O(n258));
  nor2   g0186(.a(n258), .b(n257), .O(n259));
  nor2   g0187(.a(n259), .b(n256), .O(n260));
  nor2   g0188(.a(n260), .b(n255), .O(n261));
  inv1   g0189(.a(n261), .O(n262));
  inv1   g0190(.a(G169), .O(n263));
  nor2   g0191(.a(n201), .b(n103), .O(n264));
  inv1   g0192(.a(G283), .O(n265));
  nor2   g0193(.a(n265), .b(n194), .O(n266));
  nor2   g0194(.a(n205), .b(n94), .O(n267));
  nor2   g0195(.a(n267), .b(n266), .O(n268));
  inv1   g0196(.a(n268), .O(n269));
  nor2   g0197(.a(n269), .b(n264), .O(n270));
  nor2   g0198(.a(n270), .b(n198), .O(n271));
  inv1   g0199(.a(G274), .O(n272));
  nor2   g0200(.a(n197), .b(n272), .O(n273));
  inv1   g0201(.a(n273), .O(n274));
  nor2   g0202(.a(n213), .b(G41), .O(n275));
  inv1   g0203(.a(n275), .O(n276));
  nor2   g0204(.a(n276), .b(n274), .O(n277));
  nor2   g0205(.a(n275), .b(n197), .O(n278));
  inv1   g0206(.a(n278), .O(n279));
  nor2   g0207(.a(n279), .b(n89), .O(n280));
  nor2   g0208(.a(n280), .b(n277), .O(n281));
  inv1   g0209(.a(n281), .O(n282));
  nor2   g0210(.a(n282), .b(n271), .O(n283));
  nor2   g0211(.a(n283), .b(n263), .O(n284));
  inv1   g0212(.a(G179), .O(n285));
  inv1   g0213(.a(n283), .O(n286));
  nor2   g0214(.a(n286), .b(n285), .O(n287));
  nor2   g0215(.a(n287), .b(n284), .O(n288));
  nor2   g0216(.a(n232), .b(n88), .O(n289));
  nor2   g0217(.a(n234), .b(G97), .O(n290));
  nor2   g0218(.a(n93), .b(G33), .O(n291));
  nor2   g0219(.a(n113), .b(n194), .O(n292));
  nor2   g0220(.a(n292), .b(G20), .O(n293));
  inv1   g0221(.a(n293), .O(n294));
  nor2   g0222(.a(n294), .b(n291), .O(n295));
  nor2   g0223(.a(n182), .b(n83), .O(n296));
  nor2   g0224(.a(n296), .b(n227), .O(n297));
  inv1   g0225(.a(n297), .O(n298));
  nor2   g0226(.a(n298), .b(n295), .O(n299));
  nor2   g0227(.a(n299), .b(n290), .O(n300));
  inv1   g0228(.a(n300), .O(n301));
  nor2   g0229(.a(n301), .b(n289), .O(n302));
  nor2   g0230(.a(n302), .b(n288), .O(n303));
  inv1   g0231(.a(n302), .O(n304));
  nor2   g0232(.a(n286), .b(G190), .O(n305));
  nor2   g0233(.a(n283), .b(G200), .O(n306));
  nor2   g0234(.a(n306), .b(n305), .O(n307));
  nor2   g0235(.a(n307), .b(n304), .O(n308));
  nor2   g0236(.a(n308), .b(n303), .O(n309));
  inv1   g0237(.a(n309), .O(n310));
  nor2   g0238(.a(n310), .b(n262), .O(n311));
  inv1   g0239(.a(n311), .O(n312));
  nor2   g0240(.a(n201), .b(n114), .O(n313));
  nor2   g0241(.a(n205), .b(n89), .O(n314));
  inv1   g0242(.a(G303), .O(n315));
  nor2   g0243(.a(n315), .b(n194), .O(n316));
  nor2   g0244(.a(n316), .b(n314), .O(n317));
  inv1   g0245(.a(n317), .O(n318));
  nor2   g0246(.a(n318), .b(n313), .O(n319));
  nor2   g0247(.a(n319), .b(n198), .O(n320));
  nor2   g0248(.a(n279), .b(n97), .O(n321));
  nor2   g0249(.a(n321), .b(n277), .O(n322));
  inv1   g0250(.a(n322), .O(n323));
  nor2   g0251(.a(n323), .b(n320), .O(n324));
  nor2   g0252(.a(n324), .b(G169), .O(n325));
  nor2   g0253(.a(n232), .b(n96), .O(n326));
  nor2   g0254(.a(G116), .b(n83), .O(n327));
  inv1   g0255(.a(n327), .O(n328));
  nor2   g0256(.a(n328), .b(n223), .O(n329));
  nor2   g0257(.a(n88), .b(G33), .O(n330));
  nor2   g0258(.a(n266), .b(G20), .O(n331));
  inv1   g0259(.a(n331), .O(n332));
  nor2   g0260(.a(n332), .b(n330), .O(n333));
  nor2   g0261(.a(n327), .b(n227), .O(n334));
  inv1   g0262(.a(n334), .O(n335));
  nor2   g0263(.a(n335), .b(n333), .O(n336));
  nor2   g0264(.a(n336), .b(n329), .O(n337));
  inv1   g0265(.a(n337), .O(n338));
  nor2   g0266(.a(n338), .b(n326), .O(n339));
  inv1   g0267(.a(n324), .O(n340));
  nor2   g0268(.a(n340), .b(G179), .O(n341));
  nor2   g0269(.a(n341), .b(n339), .O(n342));
  inv1   g0270(.a(n342), .O(n343));
  nor2   g0271(.a(n343), .b(n325), .O(n344));
  inv1   g0272(.a(G190), .O(n345));
  nor2   g0273(.a(n340), .b(n345), .O(n346));
  inv1   g0274(.a(n339), .O(n347));
  inv1   g0275(.a(G200), .O(n348));
  nor2   g0276(.a(n324), .b(n348), .O(n349));
  nor2   g0277(.a(n349), .b(n347), .O(n350));
  inv1   g0278(.a(n350), .O(n351));
  nor2   g0279(.a(n351), .b(n346), .O(n352));
  nor2   g0280(.a(n352), .b(n344), .O(n353));
  inv1   g0281(.a(n353), .O(n354));
  nor2   g0282(.a(n205), .b(n103), .O(n355));
  nor2   g0283(.a(n201), .b(n89), .O(n356));
  inv1   g0284(.a(G294), .O(n357));
  nor2   g0285(.a(n357), .b(n194), .O(n358));
  nor2   g0286(.a(n358), .b(n356), .O(n359));
  inv1   g0287(.a(n359), .O(n360));
  nor2   g0288(.a(n360), .b(n355), .O(n361));
  nor2   g0289(.a(n361), .b(n198), .O(n362));
  nor2   g0290(.a(n279), .b(n114), .O(n363));
  nor2   g0291(.a(n363), .b(n277), .O(n364));
  inv1   g0292(.a(n364), .O(n365));
  nor2   g0293(.a(n365), .b(n362), .O(n366));
  inv1   g0294(.a(n366), .O(n367));
  nor2   g0295(.a(n367), .b(G179), .O(n368));
  nor2   g0296(.a(n232), .b(n113), .O(n369));
  nor2   g0297(.a(n226), .b(G13), .O(n370));
  nor2   g0298(.a(G107), .b(n83), .O(n371));
  inv1   g0299(.a(n371), .O(n372));
  nor2   g0300(.a(n372), .b(n370), .O(n373));
  nor2   g0301(.a(n78), .b(G33), .O(n374));
  nor2   g0302(.a(n374), .b(n203), .O(n375));
  nor2   g0303(.a(n375), .b(G20), .O(n376));
  inv1   g0304(.a(n376), .O(n377));
  nor2   g0305(.a(n377), .b(n227), .O(n378));
  nor2   g0306(.a(n378), .b(n373), .O(n379));
  inv1   g0307(.a(n379), .O(n380));
  nor2   g0308(.a(n380), .b(n369), .O(n381));
  nor2   g0309(.a(n366), .b(G169), .O(n382));
  nor2   g0310(.a(n382), .b(n381), .O(n383));
  inv1   g0311(.a(n383), .O(n384));
  nor2   g0312(.a(n384), .b(n368), .O(n385));
  nor2   g0313(.a(n366), .b(n348), .O(n386));
  inv1   g0314(.a(n381), .O(n387));
  nor2   g0315(.a(n367), .b(n345), .O(n388));
  nor2   g0316(.a(n388), .b(n387), .O(n389));
  inv1   g0317(.a(n389), .O(n390));
  nor2   g0318(.a(n390), .b(n386), .O(n391));
  nor2   g0319(.a(n391), .b(n385), .O(n392));
  inv1   g0320(.a(n392), .O(n393));
  nor2   g0321(.a(n393), .b(n354), .O(n394));
  inv1   g0322(.a(n394), .O(n395));
  nor2   g0323(.a(n395), .b(n312), .O(n396));
  inv1   g0324(.a(n396), .O(n397));
  inv1   g0325(.a(G223), .O(n398));
  nor2   g0326(.a(n205), .b(n398), .O(n399));
  nor2   g0327(.a(n78), .b(n194), .O(n400));
  nor2   g0328(.a(n201), .b(n106), .O(n401));
  nor2   g0329(.a(n401), .b(n400), .O(n402));
  inv1   g0330(.a(n402), .O(n403));
  nor2   g0331(.a(n403), .b(n399), .O(n404));
  nor2   g0332(.a(n404), .b(n198), .O(n405));
  nor2   g0333(.a(G45), .b(G41), .O(n406));
  nor2   g0334(.a(n406), .b(G1), .O(n407));
  inv1   g0335(.a(n407), .O(n408));
  nor2   g0336(.a(n408), .b(n274), .O(n409));
  nor2   g0337(.a(n407), .b(n197), .O(n410));
  inv1   g0338(.a(n410), .O(n411));
  nor2   g0339(.a(n411), .b(n111), .O(n412));
  nor2   g0340(.a(n412), .b(n409), .O(n413));
  inv1   g0341(.a(n413), .O(n414));
  nor2   g0342(.a(n414), .b(n405), .O(n415));
  inv1   g0343(.a(n415), .O(n416));
  nor2   g0344(.a(n416), .b(G179), .O(n417));
  nor2   g0345(.a(n83), .b(G1), .O(n418));
  nor2   g0346(.a(n418), .b(n110), .O(n419));
  inv1   g0347(.a(n419), .O(n420));
  nor2   g0348(.a(n420), .b(n230), .O(n421));
  nor2   g0349(.a(n170), .b(n83), .O(n422));
  inv1   g0350(.a(G159), .O(n423));
  nor2   g0351(.a(G33), .b(G20), .O(n424));
  inv1   g0352(.a(n424), .O(n425));
  nor2   g0353(.a(n425), .b(n423), .O(n426));
  nor2   g0354(.a(n194), .b(G20), .O(n427));
  inv1   g0355(.a(n427), .O(n428));
  nor2   g0356(.a(n428), .b(n85), .O(n429));
  nor2   g0357(.a(n429), .b(n426), .O(n430));
  inv1   g0358(.a(n430), .O(n431));
  nor2   g0359(.a(n431), .b(n422), .O(n432));
  nor2   g0360(.a(n432), .b(n227), .O(n433));
  nor2   g0361(.a(n234), .b(G58), .O(n434));
  nor2   g0362(.a(n434), .b(n433), .O(n435));
  inv1   g0363(.a(n435), .O(n436));
  nor2   g0364(.a(n436), .b(n421), .O(n437));
  nor2   g0365(.a(n415), .b(G169), .O(n438));
  nor2   g0366(.a(n438), .b(n437), .O(n439));
  inv1   g0367(.a(n439), .O(n440));
  nor2   g0368(.a(n440), .b(n417), .O(n441));
  nor2   g0369(.a(n205), .b(n106), .O(n442));
  nor2   g0370(.a(n201), .b(n111), .O(n443));
  nor2   g0371(.a(n443), .b(n237), .O(n444));
  inv1   g0372(.a(n444), .O(n445));
  nor2   g0373(.a(n445), .b(n442), .O(n446));
  nor2   g0374(.a(n446), .b(n198), .O(n447));
  nor2   g0375(.a(n411), .b(n86), .O(n448));
  nor2   g0376(.a(n448), .b(n409), .O(n449));
  inv1   g0377(.a(n449), .O(n450));
  nor2   g0378(.a(n450), .b(n447), .O(n451));
  inv1   g0379(.a(n451), .O(n452));
  nor2   g0380(.a(n452), .b(G179), .O(n453));
  nor2   g0381(.a(n418), .b(n85), .O(n454));
  inv1   g0382(.a(n454), .O(n455));
  nor2   g0383(.a(n455), .b(n230), .O(n456));
  nor2   g0384(.a(n93), .b(n194), .O(n457));
  nor2   g0385(.a(n105), .b(G33), .O(n458));
  nor2   g0386(.a(n458), .b(n457), .O(n459));
  nor2   g0387(.a(n459), .b(G20), .O(n460));
  inv1   g0388(.a(n460), .O(n461));
  nor2   g0389(.a(n461), .b(n227), .O(n462));
  nor2   g0390(.a(G68), .b(n83), .O(n463));
  inv1   g0391(.a(n463), .O(n464));
  nor2   g0392(.a(n464), .b(n370), .O(n465));
  nor2   g0393(.a(n465), .b(n462), .O(n466));
  inv1   g0394(.a(n466), .O(n467));
  nor2   g0395(.a(n467), .b(n456), .O(n468));
  nor2   g0396(.a(n451), .b(G169), .O(n469));
  nor2   g0397(.a(n469), .b(n468), .O(n470));
  inv1   g0398(.a(n470), .O(n471));
  nor2   g0399(.a(n471), .b(n453), .O(n472));
  nor2   g0400(.a(n205), .b(n111), .O(n473));
  nor2   g0401(.a(n201), .b(n86), .O(n474));
  nor2   g0402(.a(n474), .b(n292), .O(n475));
  inv1   g0403(.a(n475), .O(n476));
  nor2   g0404(.a(n476), .b(n473), .O(n477));
  nor2   g0405(.a(n477), .b(n198), .O(n478));
  nor2   g0406(.a(n411), .b(n94), .O(n479));
  nor2   g0407(.a(n479), .b(n409), .O(n480));
  inv1   g0408(.a(n480), .O(n481));
  nor2   g0409(.a(n481), .b(n478), .O(n482));
  inv1   g0410(.a(n482), .O(n483));
  nor2   g0411(.a(n483), .b(G179), .O(n484));
  nor2   g0412(.a(n110), .b(G33), .O(n485));
  nor2   g0413(.a(n485), .b(G20), .O(n486));
  inv1   g0414(.a(n486), .O(n487));
  nor2   g0415(.a(n487), .b(n400), .O(n488));
  nor2   g0416(.a(G77), .b(n83), .O(n489));
  nor2   g0417(.a(n489), .b(n227), .O(n490));
  inv1   g0418(.a(n490), .O(n491));
  nor2   g0419(.a(n491), .b(n488), .O(n492));
  inv1   g0420(.a(n489), .O(n493));
  nor2   g0421(.a(n493), .b(n223), .O(n494));
  nor2   g0422(.a(n418), .b(n93), .O(n495));
  inv1   g0423(.a(n495), .O(n496));
  nor2   g0424(.a(n496), .b(n230), .O(n497));
  nor2   g0425(.a(n497), .b(n494), .O(n498));
  inv1   g0426(.a(n498), .O(n499));
  nor2   g0427(.a(n499), .b(n492), .O(n500));
  nor2   g0428(.a(n482), .b(G169), .O(n501));
  nor2   g0429(.a(n501), .b(n500), .O(n502));
  inv1   g0430(.a(n502), .O(n503));
  nor2   g0431(.a(n503), .b(n484), .O(n504));
  nor2   g0432(.a(n504), .b(n472), .O(n505));
  inv1   g0433(.a(n505), .O(n506));
  nor2   g0434(.a(n506), .b(n441), .O(n507));
  inv1   g0435(.a(n507), .O(n508));
  nor2   g0436(.a(n415), .b(n348), .O(n509));
  inv1   g0437(.a(n437), .O(n510));
  nor2   g0438(.a(n416), .b(n345), .O(n511));
  nor2   g0439(.a(n511), .b(n510), .O(n512));
  inv1   g0440(.a(n512), .O(n513));
  nor2   g0441(.a(n513), .b(n509), .O(n514));
  nor2   g0442(.a(n451), .b(n348), .O(n515));
  inv1   g0443(.a(n468), .O(n516));
  nor2   g0444(.a(n452), .b(n345), .O(n517));
  nor2   g0445(.a(n517), .b(n516), .O(n518));
  inv1   g0446(.a(n518), .O(n519));
  nor2   g0447(.a(n519), .b(n515), .O(n520));
  nor2   g0448(.a(n520), .b(n514), .O(n521));
  inv1   g0449(.a(n521), .O(n522));
  inv1   g0450(.a(G222), .O(n523));
  nor2   g0451(.a(n205), .b(n523), .O(n524));
  nor2   g0452(.a(n201), .b(n398), .O(n525));
  nor2   g0453(.a(n525), .b(n457), .O(n526));
  inv1   g0454(.a(n526), .O(n527));
  nor2   g0455(.a(n527), .b(n524), .O(n528));
  nor2   g0456(.a(n528), .b(n198), .O(n529));
  nor2   g0457(.a(n411), .b(n106), .O(n530));
  nor2   g0458(.a(n530), .b(n409), .O(n531));
  inv1   g0459(.a(n531), .O(n532));
  nor2   g0460(.a(n532), .b(n529), .O(n533));
  inv1   g0461(.a(n533), .O(n534));
  nor2   g0462(.a(n534), .b(G179), .O(n535));
  nor2   g0463(.a(n418), .b(n105), .O(n536));
  inv1   g0464(.a(n536), .O(n537));
  nor2   g0465(.a(n537), .b(n230), .O(n538));
  nor2   g0466(.a(n75), .b(n83), .O(n539));
  inv1   g0467(.a(G150), .O(n540));
  nor2   g0468(.a(n425), .b(n540), .O(n541));
  nor2   g0469(.a(n428), .b(n110), .O(n542));
  nor2   g0470(.a(n542), .b(n541), .O(n543));
  inv1   g0471(.a(n543), .O(n544));
  nor2   g0472(.a(n544), .b(n539), .O(n545));
  nor2   g0473(.a(n545), .b(n227), .O(n546));
  nor2   g0474(.a(n234), .b(G50), .O(n547));
  nor2   g0475(.a(n547), .b(n546), .O(n548));
  inv1   g0476(.a(n548), .O(n549));
  nor2   g0477(.a(n549), .b(n538), .O(n550));
  nor2   g0478(.a(n533), .b(G169), .O(n551));
  nor2   g0479(.a(n551), .b(n550), .O(n552));
  inv1   g0480(.a(n552), .O(n553));
  nor2   g0481(.a(n553), .b(n535), .O(n554));
  nor2   g0482(.a(n533), .b(n348), .O(n555));
  inv1   g0483(.a(n550), .O(n556));
  nor2   g0484(.a(n534), .b(n345), .O(n557));
  nor2   g0485(.a(n557), .b(n556), .O(n558));
  inv1   g0486(.a(n558), .O(n559));
  nor2   g0487(.a(n559), .b(n555), .O(n560));
  nor2   g0488(.a(n560), .b(n554), .O(n561));
  inv1   g0489(.a(n561), .O(n562));
  nor2   g0490(.a(n482), .b(n348), .O(n563));
  inv1   g0491(.a(n500), .O(n564));
  nor2   g0492(.a(n483), .b(n345), .O(n565));
  nor2   g0493(.a(n565), .b(n564), .O(n566));
  inv1   g0494(.a(n566), .O(n567));
  nor2   g0495(.a(n567), .b(n563), .O(n568));
  nor2   g0496(.a(n568), .b(n562), .O(n569));
  inv1   g0497(.a(n569), .O(n570));
  nor2   g0498(.a(n570), .b(n522), .O(n571));
  inv1   g0499(.a(n571), .O(n572));
  nor2   g0500(.a(n572), .b(n508), .O(n573));
  inv1   g0501(.a(n573), .O(n574));
  nor2   g0502(.a(n574), .b(n397), .O(G372));
  inv1   g0503(.a(n344), .O(n576));
  nor2   g0504(.a(n391), .b(n576), .O(n577));
  nor2   g0505(.a(n577), .b(n385), .O(n578));
  nor2   g0506(.a(n578), .b(n312), .O(n579));
  inv1   g0507(.a(n303), .O(n580));
  nor2   g0508(.a(n580), .b(n260), .O(n581));
  nor2   g0509(.a(n581), .b(n255), .O(n582));
  inv1   g0510(.a(n582), .O(n583));
  nor2   g0511(.a(n583), .b(n579), .O(n584));
  nor2   g0512(.a(n584), .b(n574), .O(n585));
  nor2   g0513(.a(n521), .b(n441), .O(n586));
  nor2   g0514(.a(n560), .b(n507), .O(n587));
  inv1   g0515(.a(n587), .O(n588));
  nor2   g0516(.a(n588), .b(n586), .O(n589));
  nor2   g0517(.a(n589), .b(n554), .O(n590));
  inv1   g0518(.a(n590), .O(n591));
  nor2   g0519(.a(n591), .b(n585), .O(n592));
  inv1   g0520(.a(n592), .O(G369));
  inv1   g0521(.a(G343), .O(n594));
  inv1   g0522(.a(G213), .O(n595));
  nor2   g0523(.a(n595), .b(G20), .O(n596));
  inv1   g0524(.a(n596), .O(n597));
  nor2   g0525(.a(n597), .b(n223), .O(n598));
  inv1   g0526(.a(n598), .O(n599));
  nor2   g0527(.a(n599), .b(n594), .O(n600));
  inv1   g0528(.a(n600), .O(n601));
  nor2   g0529(.a(n601), .b(n381), .O(n602));
  nor2   g0530(.a(n602), .b(n391), .O(n603));
  nor2   g0531(.a(n603), .b(n385), .O(n604));
  inv1   g0532(.a(G330), .O(n605));
  nor2   g0533(.a(n601), .b(n339), .O(n606));
  nor2   g0534(.a(n606), .b(n354), .O(n607));
  nor2   g0535(.a(n601), .b(n576), .O(n608));
  nor2   g0536(.a(n608), .b(n607), .O(n609));
  nor2   g0537(.a(n609), .b(n605), .O(n610));
  inv1   g0538(.a(n385), .O(n611));
  nor2   g0539(.a(n600), .b(n611), .O(n612));
  nor2   g0540(.a(n612), .b(n604), .O(n613));
  inv1   g0541(.a(n613), .O(n614));
  nor2   g0542(.a(n600), .b(n576), .O(n615));
  nor2   g0543(.a(n615), .b(n614), .O(n616));
  inv1   g0544(.a(n616), .O(n617));
  nor2   g0545(.a(n617), .b(n610), .O(n618));
  nor2   g0546(.a(n618), .b(n604), .O(G399));
  nor2   g0547(.a(n600), .b(n584), .O(n620));
  nor2   g0548(.a(n600), .b(n396), .O(n621));
  inv1   g0549(.a(n287), .O(n622));
  nor2   g0550(.a(n367), .b(n340), .O(n623));
  inv1   g0551(.a(n623), .O(n624));
  nor2   g0552(.a(n624), .b(n251), .O(n625));
  inv1   g0553(.a(n625), .O(n626));
  nor2   g0554(.a(n626), .b(n622), .O(n627));
  nor2   g0555(.a(n324), .b(G179), .O(n628));
  inv1   g0556(.a(n628), .O(n629));
  nor2   g0557(.a(n366), .b(n219), .O(n630));
  inv1   g0558(.a(n630), .O(n631));
  nor2   g0559(.a(n631), .b(n283), .O(n632));
  inv1   g0560(.a(n632), .O(n633));
  nor2   g0561(.a(n633), .b(n629), .O(n634));
  nor2   g0562(.a(n634), .b(n601), .O(n635));
  inv1   g0563(.a(n635), .O(n636));
  nor2   g0564(.a(n636), .b(n627), .O(n637));
  nor2   g0565(.a(n637), .b(n605), .O(n638));
  inv1   g0566(.a(n638), .O(n639));
  nor2   g0567(.a(n639), .b(n621), .O(n640));
  nor2   g0568(.a(n640), .b(n620), .O(n641));
  nor2   g0569(.a(n641), .b(G1), .O(n642));
  nor2   g0570(.a(n133), .b(G41), .O(n643));
  inv1   g0571(.a(n643), .O(n644));
  nor2   g0572(.a(n644), .b(n128), .O(n645));
  nor2   g0573(.a(n243), .b(G116), .O(n646));
  inv1   g0574(.a(n646), .O(n647));
  nor2   g0575(.a(n643), .b(n82), .O(n648));
  inv1   g0576(.a(n648), .O(n649));
  nor2   g0577(.a(n649), .b(n647), .O(n650));
  nor2   g0578(.a(n650), .b(n645), .O(n651));
  inv1   g0579(.a(n651), .O(n652));
  nor2   g0580(.a(n652), .b(n642), .O(n653));
  inv1   g0581(.a(n653), .O(G364));
  inv1   g0582(.a(n609), .O(n655));
  nor2   g0583(.a(n425), .b(G13), .O(n656));
  inv1   g0584(.a(n656), .O(n657));
  nor2   g0585(.a(n657), .b(n655), .O(n658));
  nor2   g0586(.a(G169), .b(n83), .O(n659));
  nor2   g0587(.a(n659), .b(n124), .O(n660));
  nor2   g0588(.a(n660), .b(n656), .O(n661));
  inv1   g0589(.a(n661), .O(n662));
  nor2   g0590(.a(n178), .b(n211), .O(n663));
  nor2   g0591(.a(n128), .b(G45), .O(n664));
  nor2   g0592(.a(n133), .b(n194), .O(n665));
  inv1   g0593(.a(n665), .O(n666));
  nor2   g0594(.a(n666), .b(n664), .O(n667));
  inv1   g0595(.a(n667), .O(n668));
  nor2   g0596(.a(n668), .b(n663), .O(n669));
  nor2   g0597(.a(n132), .b(G116), .O(n670));
  nor2   g0598(.a(n133), .b(G33), .O(n671));
  inv1   g0599(.a(n671), .O(n672));
  nor2   g0600(.a(n672), .b(n80), .O(n673));
  nor2   g0601(.a(n673), .b(n670), .O(n674));
  inv1   g0602(.a(n674), .O(n675));
  nor2   g0603(.a(n675), .b(n669), .O(n676));
  nor2   g0604(.a(n676), .b(n662), .O(n677));
  inv1   g0605(.a(n660), .O(n678));
  nor2   g0606(.a(n285), .b(n83), .O(n679));
  nor2   g0607(.a(n348), .b(n83), .O(n680));
  inv1   g0608(.a(n680), .O(n681));
  nor2   g0609(.a(n681), .b(n679), .O(n682));
  inv1   g0610(.a(n682), .O(n683));
  nor2   g0611(.a(n683), .b(n345), .O(n684));
  inv1   g0612(.a(n684), .O(n685));
  nor2   g0613(.a(n685), .b(n315), .O(n686));
  inv1   g0614(.a(G329), .O(n687));
  nor2   g0615(.a(G190), .b(n83), .O(n688));
  inv1   g0616(.a(n688), .O(n689));
  nor2   g0617(.a(n680), .b(n679), .O(n690));
  inv1   g0618(.a(n690), .O(n691));
  nor2   g0619(.a(n691), .b(n689), .O(n692));
  inv1   g0620(.a(n692), .O(n693));
  nor2   g0621(.a(n693), .b(n687), .O(n694));
  nor2   g0622(.a(n683), .b(G190), .O(n695));
  inv1   g0623(.a(n695), .O(n696));
  nor2   g0624(.a(n696), .b(n265), .O(n697));
  nor2   g0625(.a(n697), .b(n694), .O(n698));
  inv1   g0626(.a(n698), .O(n699));
  nor2   g0627(.a(n699), .b(n686), .O(n700));
  inv1   g0628(.a(n700), .O(n701));
  inv1   g0629(.a(G322), .O(n702));
  inv1   g0630(.a(n679), .O(n703));
  nor2   g0631(.a(n703), .b(G200), .O(n704));
  inv1   g0632(.a(n704), .O(n705));
  nor2   g0633(.a(n705), .b(n345), .O(n706));
  inv1   g0634(.a(n706), .O(n707));
  nor2   g0635(.a(n707), .b(n702), .O(n708));
  nor2   g0636(.a(n708), .b(n194), .O(n709));
  inv1   g0637(.a(n709), .O(n710));
  inv1   g0638(.a(G317), .O(n711));
  nor2   g0639(.a(n703), .b(n348), .O(n712));
  inv1   g0640(.a(n712), .O(n713));
  nor2   g0641(.a(n713), .b(G190), .O(n714));
  inv1   g0642(.a(n714), .O(n715));
  nor2   g0643(.a(n715), .b(n711), .O(n716));
  nor2   g0644(.a(n691), .b(n688), .O(n717));
  inv1   g0645(.a(n717), .O(n718));
  nor2   g0646(.a(n718), .b(n357), .O(n719));
  nor2   g0647(.a(n719), .b(n716), .O(n720));
  inv1   g0648(.a(n720), .O(n721));
  inv1   g0649(.a(G311), .O(n722));
  nor2   g0650(.a(n705), .b(G190), .O(n723));
  inv1   g0651(.a(n723), .O(n724));
  nor2   g0652(.a(n724), .b(n722), .O(n725));
  inv1   g0653(.a(G326), .O(n726));
  nor2   g0654(.a(n713), .b(n345), .O(n727));
  inv1   g0655(.a(n727), .O(n728));
  nor2   g0656(.a(n728), .b(n726), .O(n729));
  nor2   g0657(.a(n729), .b(n725), .O(n730));
  inv1   g0658(.a(n730), .O(n731));
  nor2   g0659(.a(n731), .b(n721), .O(n732));
  inv1   g0660(.a(n732), .O(n733));
  nor2   g0661(.a(n733), .b(n710), .O(n734));
  inv1   g0662(.a(n734), .O(n735));
  nor2   g0663(.a(n735), .b(n701), .O(n736));
  nor2   g0664(.a(n718), .b(n88), .O(n737));
  nor2   g0665(.a(n685), .b(n78), .O(n738));
  nor2   g0666(.a(n728), .b(n105), .O(n739));
  nor2   g0667(.a(n739), .b(n738), .O(n740));
  inv1   g0668(.a(n740), .O(n741));
  nor2   g0669(.a(n741), .b(n737), .O(n742));
  inv1   g0670(.a(n742), .O(n743));
  nor2   g0671(.a(n696), .b(n113), .O(n744));
  nor2   g0672(.a(n744), .b(G33), .O(n745));
  inv1   g0673(.a(n745), .O(n746));
  nor2   g0674(.a(n724), .b(n93), .O(n747));
  nor2   g0675(.a(n707), .b(n110), .O(n748));
  nor2   g0676(.a(n748), .b(n747), .O(n749));
  inv1   g0677(.a(n749), .O(n750));
  nor2   g0678(.a(n715), .b(n85), .O(n751));
  nor2   g0679(.a(n693), .b(n423), .O(n752));
  nor2   g0680(.a(n752), .b(n751), .O(n753));
  inv1   g0681(.a(n753), .O(n754));
  nor2   g0682(.a(n754), .b(n750), .O(n755));
  inv1   g0683(.a(n755), .O(n756));
  nor2   g0684(.a(n756), .b(n746), .O(n757));
  inv1   g0685(.a(n757), .O(n758));
  nor2   g0686(.a(n758), .b(n743), .O(n759));
  nor2   g0687(.a(n759), .b(n736), .O(n760));
  nor2   g0688(.a(n760), .b(n678), .O(n761));
  nor2   g0689(.a(n130), .b(n125), .O(n762));
  inv1   g0690(.a(n762), .O(n763));
  nor2   g0691(.a(n124), .b(G45), .O(n764));
  nor2   g0692(.a(n764), .b(n763), .O(n765));
  nor2   g0693(.a(n765), .b(n643), .O(n766));
  inv1   g0694(.a(n766), .O(n767));
  nor2   g0695(.a(n767), .b(n761), .O(n768));
  inv1   g0696(.a(n768), .O(n769));
  nor2   g0697(.a(n769), .b(n677), .O(n770));
  inv1   g0698(.a(n770), .O(n771));
  nor2   g0699(.a(n771), .b(n658), .O(n772));
  nor2   g0700(.a(n655), .b(G330), .O(n773));
  nor2   g0701(.a(n766), .b(n610), .O(n774));
  inv1   g0702(.a(n774), .O(n775));
  nor2   g0703(.a(n775), .b(n773), .O(n776));
  nor2   g0704(.a(n776), .b(n772), .O(n777));
  inv1   g0705(.a(n777), .O(G396));
  inv1   g0706(.a(n640), .O(n779));
  inv1   g0707(.a(n620), .O(n780));
  inv1   g0708(.a(n504), .O(n781));
  nor2   g0709(.a(n600), .b(n781), .O(n782));
  nor2   g0710(.a(n601), .b(n500), .O(n783));
  nor2   g0711(.a(n783), .b(n568), .O(n784));
  nor2   g0712(.a(n784), .b(n504), .O(n785));
  nor2   g0713(.a(n785), .b(n782), .O(n786));
  inv1   g0714(.a(n786), .O(n787));
  nor2   g0715(.a(n787), .b(n780), .O(n788));
  nor2   g0716(.a(n786), .b(n620), .O(n789));
  nor2   g0717(.a(n789), .b(n788), .O(n790));
  inv1   g0718(.a(n790), .O(n791));
  nor2   g0719(.a(n791), .b(n779), .O(n792));
  nor2   g0720(.a(n790), .b(n640), .O(n793));
  nor2   g0721(.a(n793), .b(n766), .O(n794));
  inv1   g0722(.a(n794), .O(n795));
  nor2   g0723(.a(n795), .b(n792), .O(n796));
  nor2   g0724(.a(G33), .b(G13), .O(n797));
  inv1   g0725(.a(n797), .O(n798));
  nor2   g0726(.a(n798), .b(n786), .O(n799));
  nor2   g0727(.a(n696), .b(n85), .O(n800));
  inv1   g0728(.a(G137), .O(n801));
  nor2   g0729(.a(n728), .b(n801), .O(n802));
  nor2   g0730(.a(n718), .b(n110), .O(n803));
  nor2   g0731(.a(n803), .b(n802), .O(n804));
  inv1   g0732(.a(n804), .O(n805));
  nor2   g0733(.a(n805), .b(n800), .O(n806));
  inv1   g0734(.a(n806), .O(n807));
  inv1   g0735(.a(G143), .O(n808));
  nor2   g0736(.a(n707), .b(n808), .O(n809));
  nor2   g0737(.a(n809), .b(G33), .O(n810));
  inv1   g0738(.a(n810), .O(n811));
  nor2   g0739(.a(n685), .b(n105), .O(n812));
  inv1   g0740(.a(G132), .O(n813));
  nor2   g0741(.a(n693), .b(n813), .O(n814));
  nor2   g0742(.a(n814), .b(n812), .O(n815));
  inv1   g0743(.a(n815), .O(n816));
  nor2   g0744(.a(n724), .b(n423), .O(n817));
  nor2   g0745(.a(n715), .b(n540), .O(n818));
  nor2   g0746(.a(n818), .b(n817), .O(n819));
  inv1   g0747(.a(n819), .O(n820));
  nor2   g0748(.a(n820), .b(n816), .O(n821));
  inv1   g0749(.a(n821), .O(n822));
  nor2   g0750(.a(n822), .b(n811), .O(n823));
  inv1   g0751(.a(n823), .O(n824));
  nor2   g0752(.a(n824), .b(n807), .O(n825));
  nor2   g0753(.a(n696), .b(n78), .O(n826));
  nor2   g0754(.a(n685), .b(n113), .O(n827));
  nor2   g0755(.a(n693), .b(n722), .O(n828));
  nor2   g0756(.a(n828), .b(n827), .O(n829));
  inv1   g0757(.a(n829), .O(n830));
  nor2   g0758(.a(n830), .b(n826), .O(n831));
  inv1   g0759(.a(n831), .O(n832));
  nor2   g0760(.a(n737), .b(n194), .O(n833));
  inv1   g0761(.a(n833), .O(n834));
  nor2   g0762(.a(n707), .b(n357), .O(n835));
  nor2   g0763(.a(n715), .b(n265), .O(n836));
  nor2   g0764(.a(n836), .b(n835), .O(n837));
  inv1   g0765(.a(n837), .O(n838));
  nor2   g0766(.a(n728), .b(n315), .O(n839));
  nor2   g0767(.a(n724), .b(n96), .O(n840));
  nor2   g0768(.a(n840), .b(n839), .O(n841));
  inv1   g0769(.a(n841), .O(n842));
  nor2   g0770(.a(n842), .b(n838), .O(n843));
  inv1   g0771(.a(n843), .O(n844));
  nor2   g0772(.a(n844), .b(n834), .O(n845));
  inv1   g0773(.a(n845), .O(n846));
  nor2   g0774(.a(n846), .b(n832), .O(n847));
  nor2   g0775(.a(n847), .b(n825), .O(n848));
  nor2   g0776(.a(n848), .b(n678), .O(n849));
  nor2   g0777(.a(n797), .b(n660), .O(n850));
  inv1   g0778(.a(n850), .O(n851));
  nor2   g0779(.a(n851), .b(G77), .O(n852));
  nor2   g0780(.a(n852), .b(n767), .O(n853));
  inv1   g0781(.a(n853), .O(n854));
  nor2   g0782(.a(n854), .b(n849), .O(n855));
  inv1   g0783(.a(n855), .O(n856));
  nor2   g0784(.a(n856), .b(n799), .O(n857));
  nor2   g0785(.a(n857), .b(n796), .O(n858));
  inv1   g0786(.a(n858), .O(G384));
  inv1   g0787(.a(n441), .O(n860));
  nor2   g0788(.a(n598), .b(n860), .O(n861));
  nor2   g0789(.a(n599), .b(n437), .O(n862));
  nor2   g0790(.a(n862), .b(n514), .O(n863));
  nor2   g0791(.a(n863), .b(n441), .O(n864));
  nor2   g0792(.a(n864), .b(n861), .O(n865));
  inv1   g0793(.a(n865), .O(n866));
  nor2   g0794(.a(n601), .b(n468), .O(n867));
  nor2   g0795(.a(n867), .b(n520), .O(n868));
  nor2   g0796(.a(n868), .b(n472), .O(n869));
  inv1   g0797(.a(n472), .O(n870));
  nor2   g0798(.a(n600), .b(n870), .O(n871));
  nor2   g0799(.a(n788), .b(n782), .O(n872));
  inv1   g0800(.a(n872), .O(n873));
  nor2   g0801(.a(n873), .b(n871), .O(n874));
  nor2   g0802(.a(n874), .b(n869), .O(n875));
  inv1   g0803(.a(n875), .O(n876));
  nor2   g0804(.a(n876), .b(n866), .O(n877));
  nor2   g0805(.a(n877), .b(n861), .O(n878));
  nor2   g0806(.a(n871), .b(n869), .O(n879));
  inv1   g0807(.a(n879), .O(n880));
  nor2   g0808(.a(n866), .b(n787), .O(n881));
  inv1   g0809(.a(n881), .O(n882));
  nor2   g0810(.a(n882), .b(n880), .O(n883));
  inv1   g0811(.a(n883), .O(n884));
  nor2   g0812(.a(n884), .b(n573), .O(n885));
  nor2   g0813(.a(n883), .b(n574), .O(n886));
  nor2   g0814(.a(n886), .b(n885), .O(n887));
  nor2   g0815(.a(n887), .b(n779), .O(n888));
  inv1   g0816(.a(n888), .O(n889));
  nor2   g0817(.a(n889), .b(n878), .O(n890));
  inv1   g0818(.a(n878), .O(n891));
  nor2   g0819(.a(n888), .b(n891), .O(n892));
  nor2   g0820(.a(n892), .b(n890), .O(n893));
  nor2   g0821(.a(n780), .b(n574), .O(n894));
  nor2   g0822(.a(n894), .b(n591), .O(n895));
  inv1   g0823(.a(n895), .O(n896));
  nor2   g0824(.a(n896), .b(n893), .O(n897));
  inv1   g0825(.a(n893), .O(n898));
  nor2   g0826(.a(n895), .b(n898), .O(n899));
  nor2   g0827(.a(n899), .b(n763), .O(n900));
  inv1   g0828(.a(n900), .O(n901));
  nor2   g0829(.a(n901), .b(n897), .O(n902));
  nor2   g0830(.a(n172), .b(n105), .O(n903));
  nor2   g0831(.a(G68), .b(G50), .O(n904));
  nor2   g0832(.a(n904), .b(n131), .O(n905));
  inv1   g0833(.a(n905), .O(n906));
  nor2   g0834(.a(n906), .b(n903), .O(n907));
  inv1   g0835(.a(n296), .O(n908));
  nor2   g0836(.a(n124), .b(n96), .O(n909));
  inv1   g0837(.a(n909), .O(n910));
  nor2   g0838(.a(n910), .b(n908), .O(n911));
  nor2   g0839(.a(n911), .b(n907), .O(n912));
  inv1   g0840(.a(n912), .O(n913));
  nor2   g0841(.a(n913), .b(n902), .O(n914));
  inv1   g0842(.a(n914), .O(G367));
  nor2   g0843(.a(n601), .b(n250), .O(n916));
  nor2   g0844(.a(n916), .b(n262), .O(n917));
  inv1   g0845(.a(n255), .O(n918));
  nor2   g0846(.a(n601), .b(n918), .O(n919));
  nor2   g0847(.a(n919), .b(n917), .O(n920));
  inv1   g0848(.a(n920), .O(n921));
  nor2   g0849(.a(n921), .b(n657), .O(n922));
  nor2   g0850(.a(n696), .b(n88), .O(n923));
  nor2   g0851(.a(n715), .b(n357), .O(n924));
  nor2   g0852(.a(n718), .b(n113), .O(n925));
  nor2   g0853(.a(n925), .b(n924), .O(n926));
  inv1   g0854(.a(n926), .O(n927));
  nor2   g0855(.a(n927), .b(n923), .O(n928));
  inv1   g0856(.a(n928), .O(n929));
  nor2   g0857(.a(n707), .b(n315), .O(n930));
  nor2   g0858(.a(n930), .b(n194), .O(n931));
  inv1   g0859(.a(n931), .O(n932));
  nor2   g0860(.a(n685), .b(n96), .O(n933));
  nor2   g0861(.a(n728), .b(n722), .O(n934));
  nor2   g0862(.a(n934), .b(n933), .O(n935));
  inv1   g0863(.a(n935), .O(n936));
  nor2   g0864(.a(n693), .b(n711), .O(n937));
  nor2   g0865(.a(n724), .b(n265), .O(n938));
  nor2   g0866(.a(n938), .b(n937), .O(n939));
  inv1   g0867(.a(n939), .O(n940));
  nor2   g0868(.a(n940), .b(n936), .O(n941));
  inv1   g0869(.a(n941), .O(n942));
  nor2   g0870(.a(n942), .b(n932), .O(n943));
  inv1   g0871(.a(n943), .O(n944));
  nor2   g0872(.a(n944), .b(n929), .O(n945));
  nor2   g0873(.a(n724), .b(n105), .O(n946));
  nor2   g0874(.a(n715), .b(n423), .O(n947));
  nor2   g0875(.a(n728), .b(n808), .O(n948));
  nor2   g0876(.a(n948), .b(n947), .O(n949));
  inv1   g0877(.a(n949), .O(n950));
  nor2   g0878(.a(n950), .b(n946), .O(n951));
  inv1   g0879(.a(n951), .O(n952));
  nor2   g0880(.a(n696), .b(n93), .O(n953));
  nor2   g0881(.a(n953), .b(G33), .O(n954));
  inv1   g0882(.a(n954), .O(n955));
  nor2   g0883(.a(n693), .b(n801), .O(n956));
  nor2   g0884(.a(n718), .b(n85), .O(n957));
  nor2   g0885(.a(n957), .b(n956), .O(n958));
  inv1   g0886(.a(n958), .O(n959));
  nor2   g0887(.a(n707), .b(n540), .O(n960));
  nor2   g0888(.a(n685), .b(n110), .O(n961));
  nor2   g0889(.a(n961), .b(n960), .O(n962));
  inv1   g0890(.a(n962), .O(n963));
  nor2   g0891(.a(n963), .b(n959), .O(n964));
  inv1   g0892(.a(n964), .O(n965));
  nor2   g0893(.a(n965), .b(n955), .O(n966));
  inv1   g0894(.a(n966), .O(n967));
  nor2   g0895(.a(n967), .b(n952), .O(n968));
  nor2   g0896(.a(n968), .b(n945), .O(n969));
  nor2   g0897(.a(n969), .b(n678), .O(n970));
  nor2   g0898(.a(n666), .b(n151), .O(n971));
  nor2   g0899(.a(n132), .b(n78), .O(n972));
  nor2   g0900(.a(n972), .b(n662), .O(n973));
  inv1   g0901(.a(n973), .O(n974));
  nor2   g0902(.a(n974), .b(n971), .O(n975));
  nor2   g0903(.a(n975), .b(n767), .O(n976));
  inv1   g0904(.a(n976), .O(n977));
  nor2   g0905(.a(n977), .b(n970), .O(n978));
  inv1   g0906(.a(n978), .O(n979));
  nor2   g0907(.a(n979), .b(n922), .O(n980));
  inv1   g0908(.a(n641), .O(n981));
  inv1   g0909(.a(n610), .O(n982));
  inv1   g0910(.a(n615), .O(n983));
  nor2   g0911(.a(n983), .b(n613), .O(n984));
  nor2   g0912(.a(n984), .b(n616), .O(n985));
  inv1   g0913(.a(n985), .O(n986));
  nor2   g0914(.a(n986), .b(n982), .O(n987));
  nor2   g0915(.a(n985), .b(n610), .O(n988));
  nor2   g0916(.a(n988), .b(n987), .O(n989));
  nor2   g0917(.a(n989), .b(n981), .O(n990));
  inv1   g0918(.a(n990), .O(n991));
  nor2   g0919(.a(n600), .b(n580), .O(n992));
  nor2   g0920(.a(n601), .b(n302), .O(n993));
  nor2   g0921(.a(n993), .b(n308), .O(n994));
  nor2   g0922(.a(n994), .b(n303), .O(n995));
  nor2   g0923(.a(n995), .b(n992), .O(n996));
  inv1   g0924(.a(n996), .O(n997));
  nor2   g0925(.a(n997), .b(G399), .O(n998));
  inv1   g0926(.a(G399), .O(n999));
  nor2   g0927(.a(n996), .b(n999), .O(n1000));
  nor2   g0928(.a(n1000), .b(n998), .O(n1001));
  nor2   g0929(.a(n1001), .b(n991), .O(n1002));
  nor2   g0930(.a(n765), .b(n981), .O(n1003));
  inv1   g0931(.a(n1003), .O(n1004));
  nor2   g0932(.a(n1004), .b(n1002), .O(n1005));
  nor2   g0933(.a(n998), .b(n995), .O(n1006));
  nor2   g0934(.a(n1006), .b(n921), .O(n1007));
  inv1   g0935(.a(n1006), .O(n1008));
  nor2   g0936(.a(n1008), .b(n920), .O(n1009));
  nor2   g0937(.a(n1009), .b(n766), .O(n1010));
  inv1   g0938(.a(n1010), .O(n1011));
  nor2   g0939(.a(n1011), .b(n1007), .O(n1012));
  inv1   g0940(.a(n1012), .O(n1013));
  nor2   g0941(.a(n1013), .b(n1005), .O(n1014));
  nor2   g0942(.a(n1014), .b(n980), .O(n1015));
  inv1   g0943(.a(n1015), .O(G387));
  inv1   g0944(.a(n989), .O(n1017));
  nor2   g0945(.a(n1017), .b(n641), .O(n1018));
  nor2   g0946(.a(n990), .b(n644), .O(n1019));
  inv1   g0947(.a(n1019), .O(n1020));
  nor2   g0948(.a(n1020), .b(n1018), .O(n1021));
  inv1   g0949(.a(n765), .O(n1022));
  nor2   g0950(.a(n989), .b(n1022), .O(n1023));
  nor2   g0951(.a(n657), .b(n613), .O(n1024));
  nor2   g0952(.a(n707), .b(n105), .O(n1025));
  nor2   g0953(.a(n724), .b(n85), .O(n1026));
  nor2   g0954(.a(n685), .b(n93), .O(n1027));
  nor2   g0955(.a(n1027), .b(n1026), .O(n1028));
  inv1   g0956(.a(n1028), .O(n1029));
  nor2   g0957(.a(n1029), .b(n1025), .O(n1030));
  inv1   g0958(.a(n1030), .O(n1031));
  nor2   g0959(.a(n923), .b(G33), .O(n1032));
  inv1   g0960(.a(n1032), .O(n1033));
  nor2   g0961(.a(n715), .b(n110), .O(n1034));
  nor2   g0962(.a(n693), .b(n540), .O(n1035));
  nor2   g0963(.a(n1035), .b(n1034), .O(n1036));
  inv1   g0964(.a(n1036), .O(n1037));
  nor2   g0965(.a(n728), .b(n423), .O(n1038));
  nor2   g0966(.a(n718), .b(n78), .O(n1039));
  nor2   g0967(.a(n1039), .b(n1038), .O(n1040));
  inv1   g0968(.a(n1040), .O(n1041));
  nor2   g0969(.a(n1041), .b(n1037), .O(n1042));
  inv1   g0970(.a(n1042), .O(n1043));
  nor2   g0971(.a(n1043), .b(n1033), .O(n1044));
  inv1   g0972(.a(n1044), .O(n1045));
  nor2   g0973(.a(n1045), .b(n1031), .O(n1046));
  nor2   g0974(.a(n685), .b(n357), .O(n1047));
  nor2   g0975(.a(n728), .b(n702), .O(n1048));
  nor2   g0976(.a(n718), .b(n265), .O(n1049));
  nor2   g0977(.a(n1049), .b(n1048), .O(n1050));
  inv1   g0978(.a(n1050), .O(n1051));
  nor2   g0979(.a(n1051), .b(n1047), .O(n1052));
  inv1   g0980(.a(n1052), .O(n1053));
  nor2   g0981(.a(n707), .b(n711), .O(n1054));
  nor2   g0982(.a(n1054), .b(n194), .O(n1055));
  inv1   g0983(.a(n1055), .O(n1056));
  nor2   g0984(.a(n715), .b(n722), .O(n1057));
  nor2   g0985(.a(n696), .b(n96), .O(n1058));
  nor2   g0986(.a(n1058), .b(n1057), .O(n1059));
  inv1   g0987(.a(n1059), .O(n1060));
  nor2   g0988(.a(n693), .b(n726), .O(n1061));
  nor2   g0989(.a(n724), .b(n315), .O(n1062));
  nor2   g0990(.a(n1062), .b(n1061), .O(n1063));
  inv1   g0991(.a(n1063), .O(n1064));
  nor2   g0992(.a(n1064), .b(n1060), .O(n1065));
  inv1   g0993(.a(n1065), .O(n1066));
  nor2   g0994(.a(n1066), .b(n1056), .O(n1067));
  inv1   g0995(.a(n1067), .O(n1068));
  nor2   g0996(.a(n1068), .b(n1053), .O(n1069));
  nor2   g0997(.a(n1069), .b(n1046), .O(n1070));
  nor2   g0998(.a(n1070), .b(n678), .O(n1071));
  nor2   g0999(.a(n163), .b(n211), .O(n1072));
  nor2   g1000(.a(n93), .b(n85), .O(n1073));
  nor2   g1001(.a(G50), .b(G45), .O(n1074));
  inv1   g1002(.a(n1074), .O(n1075));
  nor2   g1003(.a(n1075), .b(n110), .O(n1076));
  inv1   g1004(.a(n1076), .O(n1077));
  nor2   g1005(.a(n1077), .b(n1073), .O(n1078));
  inv1   g1006(.a(n1078), .O(n1079));
  nor2   g1007(.a(n1079), .b(n647), .O(n1080));
  nor2   g1008(.a(n1080), .b(n666), .O(n1081));
  inv1   g1009(.a(n1081), .O(n1082));
  nor2   g1010(.a(n1082), .b(n1072), .O(n1083));
  nor2   g1011(.a(n132), .b(G107), .O(n1084));
  nor2   g1012(.a(n672), .b(n646), .O(n1085));
  nor2   g1013(.a(n1085), .b(n1084), .O(n1086));
  inv1   g1014(.a(n1086), .O(n1087));
  nor2   g1015(.a(n1087), .b(n1083), .O(n1088));
  nor2   g1016(.a(n1088), .b(n662), .O(n1089));
  nor2   g1017(.a(n1089), .b(n767), .O(n1090));
  inv1   g1018(.a(n1090), .O(n1091));
  nor2   g1019(.a(n1091), .b(n1071), .O(n1092));
  inv1   g1020(.a(n1092), .O(n1093));
  nor2   g1021(.a(n1093), .b(n1024), .O(n1094));
  nor2   g1022(.a(n1094), .b(n1023), .O(n1095));
  inv1   g1023(.a(n1095), .O(n1096));
  nor2   g1024(.a(n1096), .b(n1021), .O(n1097));
  inv1   g1025(.a(n1097), .O(G393));
  inv1   g1026(.a(n1001), .O(n1099));
  nor2   g1027(.a(n1099), .b(n990), .O(n1100));
  nor2   g1028(.a(n1002), .b(n644), .O(n1101));
  inv1   g1029(.a(n1101), .O(n1102));
  nor2   g1030(.a(n1102), .b(n1100), .O(n1103));
  nor2   g1031(.a(n1001), .b(n1022), .O(n1104));
  nor2   g1032(.a(n996), .b(n657), .O(n1105));
  nor2   g1033(.a(n728), .b(n540), .O(n1106));
  nor2   g1034(.a(n693), .b(n808), .O(n1107));
  nor2   g1035(.a(n707), .b(n423), .O(n1108));
  nor2   g1036(.a(n1108), .b(n1107), .O(n1109));
  inv1   g1037(.a(n1109), .O(n1110));
  nor2   g1038(.a(n1110), .b(n1106), .O(n1111));
  inv1   g1039(.a(n1111), .O(n1112));
  nor2   g1040(.a(n826), .b(G33), .O(n1113));
  inv1   g1041(.a(n1113), .O(n1114));
  nor2   g1042(.a(n685), .b(n85), .O(n1115));
  nor2   g1043(.a(n724), .b(n110), .O(n1116));
  nor2   g1044(.a(n1116), .b(n1115), .O(n1117));
  inv1   g1045(.a(n1117), .O(n1118));
  nor2   g1046(.a(n718), .b(n93), .O(n1119));
  nor2   g1047(.a(n715), .b(n105), .O(n1120));
  nor2   g1048(.a(n1120), .b(n1119), .O(n1121));
  inv1   g1049(.a(n1121), .O(n1122));
  nor2   g1050(.a(n1122), .b(n1118), .O(n1123));
  inv1   g1051(.a(n1123), .O(n1124));
  nor2   g1052(.a(n1124), .b(n1114), .O(n1125));
  inv1   g1053(.a(n1125), .O(n1126));
  nor2   g1054(.a(n1126), .b(n1112), .O(n1127));
  nor2   g1055(.a(n728), .b(n711), .O(n1128));
  nor2   g1056(.a(n693), .b(n702), .O(n1129));
  nor2   g1057(.a(n707), .b(n722), .O(n1130));
  nor2   g1058(.a(n1130), .b(n1129), .O(n1131));
  inv1   g1059(.a(n1131), .O(n1132));
  nor2   g1060(.a(n1132), .b(n1128), .O(n1133));
  inv1   g1061(.a(n1133), .O(n1134));
  nor2   g1062(.a(n744), .b(n194), .O(n1135));
  inv1   g1063(.a(n1135), .O(n1136));
  nor2   g1064(.a(n685), .b(n265), .O(n1137));
  nor2   g1065(.a(n724), .b(n357), .O(n1138));
  nor2   g1066(.a(n1138), .b(n1137), .O(n1139));
  inv1   g1067(.a(n1139), .O(n1140));
  nor2   g1068(.a(n718), .b(n96), .O(n1141));
  nor2   g1069(.a(n715), .b(n315), .O(n1142));
  nor2   g1070(.a(n1142), .b(n1141), .O(n1143));
  inv1   g1071(.a(n1143), .O(n1144));
  nor2   g1072(.a(n1144), .b(n1140), .O(n1145));
  inv1   g1073(.a(n1145), .O(n1146));
  nor2   g1074(.a(n1146), .b(n1136), .O(n1147));
  inv1   g1075(.a(n1147), .O(n1148));
  nor2   g1076(.a(n1148), .b(n1134), .O(n1149));
  nor2   g1077(.a(n1149), .b(n1127), .O(n1150));
  nor2   g1078(.a(n1150), .b(n678), .O(n1151));
  nor2   g1079(.a(n666), .b(n190), .O(n1152));
  nor2   g1080(.a(n132), .b(n88), .O(n1153));
  nor2   g1081(.a(n1153), .b(n662), .O(n1154));
  inv1   g1082(.a(n1154), .O(n1155));
  nor2   g1083(.a(n1155), .b(n1152), .O(n1156));
  nor2   g1084(.a(n1156), .b(n767), .O(n1157));
  inv1   g1085(.a(n1157), .O(n1158));
  nor2   g1086(.a(n1158), .b(n1151), .O(n1159));
  inv1   g1087(.a(n1159), .O(n1160));
  nor2   g1088(.a(n1160), .b(n1105), .O(n1161));
  nor2   g1089(.a(n1161), .b(n1104), .O(n1162));
  inv1   g1090(.a(n1162), .O(n1163));
  nor2   g1091(.a(n1163), .b(n1103), .O(n1164));
  inv1   g1092(.a(n1164), .O(G390));
  nor2   g1093(.a(n875), .b(n865), .O(n1166));
  nor2   g1094(.a(n1166), .b(n877), .O(n1167));
  nor2   g1095(.a(n787), .b(n779), .O(n1168));
  inv1   g1096(.a(n1168), .O(n1169));
  nor2   g1097(.a(n1169), .b(n880), .O(n1170));
  inv1   g1098(.a(n1170), .O(n1171));
  nor2   g1099(.a(n1171), .b(n1167), .O(n1172));
  inv1   g1100(.a(n1167), .O(n1173));
  nor2   g1101(.a(n1170), .b(n1173), .O(n1174));
  nor2   g1102(.a(n1174), .b(n1172), .O(n1175));
  inv1   g1103(.a(n1175), .O(n1176));
  nor2   g1104(.a(n641), .b(n574), .O(n1177));
  nor2   g1105(.a(n1177), .b(n591), .O(n1178));
  inv1   g1106(.a(n1178), .O(n1179));
  nor2   g1107(.a(n1168), .b(n879), .O(n1180));
  nor2   g1108(.a(n1180), .b(n1170), .O(n1181));
  nor2   g1109(.a(n1181), .b(n873), .O(n1182));
  inv1   g1110(.a(n1181), .O(n1183));
  nor2   g1111(.a(n1183), .b(n872), .O(n1184));
  nor2   g1112(.a(n1184), .b(n1182), .O(n1185));
  inv1   g1113(.a(n1185), .O(n1186));
  nor2   g1114(.a(n1186), .b(n1179), .O(n1187));
  nor2   g1115(.a(n1187), .b(n1176), .O(n1188));
  inv1   g1116(.a(n1187), .O(n1189));
  nor2   g1117(.a(n1189), .b(n1175), .O(n1190));
  nor2   g1118(.a(n1190), .b(n644), .O(n1191));
  inv1   g1119(.a(n1191), .O(n1192));
  nor2   g1120(.a(n1192), .b(n1188), .O(n1193));
  nor2   g1121(.a(n1175), .b(n1022), .O(n1194));
  nor2   g1122(.a(n865), .b(n798), .O(n1195));
  nor2   g1123(.a(n696), .b(n105), .O(n1196));
  inv1   g1124(.a(G128), .O(n1197));
  nor2   g1125(.a(n728), .b(n1197), .O(n1198));
  nor2   g1126(.a(n718), .b(n423), .O(n1199));
  nor2   g1127(.a(n1199), .b(n1198), .O(n1200));
  inv1   g1128(.a(n1200), .O(n1201));
  nor2   g1129(.a(n1201), .b(n1196), .O(n1202));
  inv1   g1130(.a(n1202), .O(n1203));
  nor2   g1131(.a(n707), .b(n813), .O(n1204));
  nor2   g1132(.a(n1204), .b(G33), .O(n1205));
  inv1   g1133(.a(n1205), .O(n1206));
  nor2   g1134(.a(n685), .b(n540), .O(n1207));
  inv1   g1135(.a(G125), .O(n1208));
  nor2   g1136(.a(n693), .b(n1208), .O(n1209));
  nor2   g1137(.a(n1209), .b(n1207), .O(n1210));
  inv1   g1138(.a(n1210), .O(n1211));
  nor2   g1139(.a(n724), .b(n808), .O(n1212));
  nor2   g1140(.a(n715), .b(n801), .O(n1213));
  nor2   g1141(.a(n1213), .b(n1212), .O(n1214));
  inv1   g1142(.a(n1214), .O(n1215));
  nor2   g1143(.a(n1215), .b(n1211), .O(n1216));
  inv1   g1144(.a(n1216), .O(n1217));
  nor2   g1145(.a(n1217), .b(n1206), .O(n1218));
  inv1   g1146(.a(n1218), .O(n1219));
  nor2   g1147(.a(n1219), .b(n1203), .O(n1220));
  nor2   g1148(.a(n707), .b(n96), .O(n1221));
  nor2   g1149(.a(n693), .b(n357), .O(n1222));
  nor2   g1150(.a(n724), .b(n88), .O(n1223));
  nor2   g1151(.a(n1223), .b(n1222), .O(n1224));
  inv1   g1152(.a(n1224), .O(n1225));
  nor2   g1153(.a(n1225), .b(n1221), .O(n1226));
  inv1   g1154(.a(n1226), .O(n1227));
  nor2   g1155(.a(n738), .b(n194), .O(n1228));
  inv1   g1156(.a(n1228), .O(n1229));
  nor2   g1157(.a(n1119), .b(n800), .O(n1230));
  inv1   g1158(.a(n1230), .O(n1231));
  nor2   g1159(.a(n715), .b(n113), .O(n1232));
  nor2   g1160(.a(n728), .b(n265), .O(n1233));
  nor2   g1161(.a(n1233), .b(n1232), .O(n1234));
  inv1   g1162(.a(n1234), .O(n1235));
  nor2   g1163(.a(n1235), .b(n1231), .O(n1236));
  inv1   g1164(.a(n1236), .O(n1237));
  nor2   g1165(.a(n1237), .b(n1229), .O(n1238));
  inv1   g1166(.a(n1238), .O(n1239));
  nor2   g1167(.a(n1239), .b(n1227), .O(n1240));
  nor2   g1168(.a(n1240), .b(n1220), .O(n1241));
  nor2   g1169(.a(n1241), .b(n678), .O(n1242));
  nor2   g1170(.a(n851), .b(G58), .O(n1243));
  nor2   g1171(.a(n1243), .b(n767), .O(n1244));
  inv1   g1172(.a(n1244), .O(n1245));
  nor2   g1173(.a(n1245), .b(n1242), .O(n1246));
  inv1   g1174(.a(n1246), .O(n1247));
  nor2   g1175(.a(n1247), .b(n1195), .O(n1248));
  nor2   g1176(.a(n1248), .b(n1194), .O(n1249));
  inv1   g1177(.a(n1249), .O(n1250));
  nor2   g1178(.a(n1250), .b(n1193), .O(n1251));
  inv1   g1179(.a(n1251), .O(G378));
  nor2   g1180(.a(n1190), .b(n1179), .O(n1253));
  nor2   g1181(.a(n599), .b(n550), .O(n1254));
  nor2   g1182(.a(n1254), .b(n562), .O(n1255));
  inv1   g1183(.a(n554), .O(n1256));
  nor2   g1184(.a(n599), .b(n1256), .O(n1257));
  nor2   g1185(.a(n1257), .b(n1255), .O(n1258));
  inv1   g1186(.a(n1258), .O(n1259));
  nor2   g1187(.a(n884), .b(n779), .O(n1260));
  nor2   g1188(.a(n1260), .b(n891), .O(n1261));
  inv1   g1189(.a(n877), .O(n1262));
  nor2   g1190(.a(n1171), .b(n1262), .O(n1263));
  nor2   g1191(.a(n1263), .b(n1261), .O(n1264));
  inv1   g1192(.a(n1264), .O(n1265));
  nor2   g1193(.a(n1265), .b(n1259), .O(n1266));
  nor2   g1194(.a(n1264), .b(n1258), .O(n1267));
  nor2   g1195(.a(n1267), .b(n1266), .O(n1268));
  nor2   g1196(.a(n1268), .b(n644), .O(n1269));
  inv1   g1197(.a(n1269), .O(n1270));
  nor2   g1198(.a(n1270), .b(n1253), .O(n1271));
  nor2   g1199(.a(n1268), .b(n1022), .O(n1272));
  nor2   g1200(.a(n1259), .b(n798), .O(n1273));
  nor2   g1201(.a(n724), .b(n801), .O(n1274));
  inv1   g1202(.a(G124), .O(n1275));
  nor2   g1203(.a(n693), .b(n1275), .O(n1276));
  nor2   g1204(.a(n696), .b(n423), .O(n1277));
  nor2   g1205(.a(n1277), .b(n1276), .O(n1278));
  inv1   g1206(.a(n1278), .O(n1279));
  nor2   g1207(.a(n1279), .b(n1274), .O(n1280));
  inv1   g1208(.a(n1280), .O(n1281));
  nor2   g1209(.a(n718), .b(n540), .O(n1282));
  nor2   g1210(.a(G41), .b(G33), .O(n1283));
  inv1   g1211(.a(n1283), .O(n1284));
  nor2   g1212(.a(n1284), .b(n1282), .O(n1285));
  inv1   g1213(.a(n1285), .O(n1286));
  nor2   g1214(.a(n685), .b(n808), .O(n1287));
  nor2   g1215(.a(n707), .b(n1197), .O(n1288));
  nor2   g1216(.a(n1288), .b(n1287), .O(n1289));
  inv1   g1217(.a(n1289), .O(n1290));
  nor2   g1218(.a(n715), .b(n813), .O(n1291));
  nor2   g1219(.a(n728), .b(n1208), .O(n1292));
  nor2   g1220(.a(n1292), .b(n1291), .O(n1293));
  inv1   g1221(.a(n1293), .O(n1294));
  nor2   g1222(.a(n1294), .b(n1290), .O(n1295));
  inv1   g1223(.a(n1295), .O(n1296));
  nor2   g1224(.a(n1296), .b(n1286), .O(n1297));
  inv1   g1225(.a(n1297), .O(n1298));
  nor2   g1226(.a(n1298), .b(n1281), .O(n1299));
  nor2   g1227(.a(G50), .b(n195), .O(n1300));
  nor2   g1228(.a(n707), .b(n113), .O(n1301));
  nor2   g1229(.a(n724), .b(n78), .O(n1302));
  nor2   g1230(.a(n693), .b(n265), .O(n1303));
  nor2   g1231(.a(n1303), .b(n1302), .O(n1304));
  inv1   g1232(.a(n1304), .O(n1305));
  nor2   g1233(.a(n1305), .b(n1301), .O(n1306));
  inv1   g1234(.a(n1306), .O(n1307));
  nor2   g1235(.a(G41), .b(n194), .O(n1308));
  inv1   g1236(.a(n1308), .O(n1309));
  nor2   g1237(.a(n1309), .b(n957), .O(n1310));
  inv1   g1238(.a(n1310), .O(n1311));
  nor2   g1239(.a(n715), .b(n88), .O(n1312));
  nor2   g1240(.a(n1312), .b(n1027), .O(n1313));
  inv1   g1241(.a(n1313), .O(n1314));
  nor2   g1242(.a(n696), .b(n110), .O(n1315));
  nor2   g1243(.a(n728), .b(n96), .O(n1316));
  nor2   g1244(.a(n1316), .b(n1315), .O(n1317));
  inv1   g1245(.a(n1317), .O(n1318));
  nor2   g1246(.a(n1318), .b(n1314), .O(n1319));
  inv1   g1247(.a(n1319), .O(n1320));
  nor2   g1248(.a(n1320), .b(n1311), .O(n1321));
  inv1   g1249(.a(n1321), .O(n1322));
  nor2   g1250(.a(n1322), .b(n1307), .O(n1323));
  nor2   g1251(.a(n1323), .b(n1300), .O(n1324));
  inv1   g1252(.a(n1324), .O(n1325));
  nor2   g1253(.a(n1325), .b(n1299), .O(n1326));
  nor2   g1254(.a(n1326), .b(n678), .O(n1327));
  nor2   g1255(.a(n851), .b(G50), .O(n1328));
  nor2   g1256(.a(n1328), .b(n767), .O(n1329));
  inv1   g1257(.a(n1329), .O(n1330));
  nor2   g1258(.a(n1330), .b(n1327), .O(n1331));
  inv1   g1259(.a(n1331), .O(n1332));
  nor2   g1260(.a(n1332), .b(n1273), .O(n1333));
  nor2   g1261(.a(n1333), .b(n1272), .O(n1334));
  inv1   g1262(.a(n1334), .O(n1335));
  nor2   g1263(.a(n1335), .b(n1271), .O(n1336));
  inv1   g1264(.a(n1336), .O(G375));
  nor2   g1265(.a(n1185), .b(n1178), .O(n1338));
  nor2   g1266(.a(n1187), .b(n644), .O(n1339));
  inv1   g1267(.a(n1339), .O(n1340));
  nor2   g1268(.a(n1340), .b(n1338), .O(n1341));
  nor2   g1269(.a(n1186), .b(n1022), .O(n1342));
  nor2   g1270(.a(n879), .b(n798), .O(n1343));
  nor2   g1271(.a(n718), .b(n105), .O(n1344));
  nor2   g1272(.a(n707), .b(n801), .O(n1345));
  nor2   g1273(.a(n724), .b(n540), .O(n1346));
  nor2   g1274(.a(n1346), .b(n1345), .O(n1347));
  inv1   g1275(.a(n1347), .O(n1348));
  nor2   g1276(.a(n1348), .b(n1344), .O(n1349));
  inv1   g1277(.a(n1349), .O(n1350));
  nor2   g1278(.a(n1315), .b(G33), .O(n1351));
  inv1   g1279(.a(n1351), .O(n1352));
  nor2   g1280(.a(n685), .b(n423), .O(n1353));
  nor2   g1281(.a(n693), .b(n1197), .O(n1354));
  nor2   g1282(.a(n1354), .b(n1353), .O(n1355));
  inv1   g1283(.a(n1355), .O(n1356));
  nor2   g1284(.a(n715), .b(n808), .O(n1357));
  nor2   g1285(.a(n728), .b(n813), .O(n1358));
  nor2   g1286(.a(n1358), .b(n1357), .O(n1359));
  inv1   g1287(.a(n1359), .O(n1360));
  nor2   g1288(.a(n1360), .b(n1356), .O(n1361));
  inv1   g1289(.a(n1361), .O(n1362));
  nor2   g1290(.a(n1362), .b(n1352), .O(n1363));
  inv1   g1291(.a(n1363), .O(n1364));
  nor2   g1292(.a(n1364), .b(n1350), .O(n1365));
  nor2   g1293(.a(n707), .b(n265), .O(n1366));
  nor2   g1294(.a(n728), .b(n357), .O(n1367));
  nor2   g1295(.a(n715), .b(n96), .O(n1368));
  nor2   g1296(.a(n1368), .b(n1367), .O(n1369));
  inv1   g1297(.a(n1369), .O(n1370));
  nor2   g1298(.a(n1370), .b(n1366), .O(n1371));
  inv1   g1299(.a(n1371), .O(n1372));
  nor2   g1300(.a(n953), .b(n194), .O(n1373));
  inv1   g1301(.a(n1373), .O(n1374));
  nor2   g1302(.a(n685), .b(n88), .O(n1375));
  nor2   g1303(.a(n1375), .b(n1039), .O(n1376));
  inv1   g1304(.a(n1376), .O(n1377));
  nor2   g1305(.a(n693), .b(n315), .O(n1378));
  nor2   g1306(.a(n724), .b(n113), .O(n1379));
  nor2   g1307(.a(n1379), .b(n1378), .O(n1380));
  inv1   g1308(.a(n1380), .O(n1381));
  nor2   g1309(.a(n1381), .b(n1377), .O(n1382));
  inv1   g1310(.a(n1382), .O(n1383));
  nor2   g1311(.a(n1383), .b(n1374), .O(n1384));
  inv1   g1312(.a(n1384), .O(n1385));
  nor2   g1313(.a(n1385), .b(n1372), .O(n1386));
  nor2   g1314(.a(n1386), .b(n1365), .O(n1387));
  nor2   g1315(.a(n1387), .b(n678), .O(n1388));
  nor2   g1316(.a(n851), .b(G68), .O(n1389));
  nor2   g1317(.a(n1389), .b(n767), .O(n1390));
  inv1   g1318(.a(n1390), .O(n1391));
  nor2   g1319(.a(n1391), .b(n1388), .O(n1392));
  inv1   g1320(.a(n1392), .O(n1393));
  nor2   g1321(.a(n1393), .b(n1343), .O(n1394));
  nor2   g1322(.a(n1394), .b(n1342), .O(n1395));
  inv1   g1323(.a(n1395), .O(n1396));
  nor2   g1324(.a(n1396), .b(n1341), .O(n1397));
  inv1   g1325(.a(n1397), .O(G381));
  nor2   g1326(.a(G375), .b(G378), .O(n1399));
  inv1   g1327(.a(n1399), .O(n1400));
  nor2   g1328(.a(G381), .b(G384), .O(n1401));
  inv1   g1329(.a(n1401), .O(n1402));
  nor2   g1330(.a(G390), .b(G387), .O(n1403));
  inv1   g1331(.a(n1403), .O(n1404));
  nor2   g1332(.a(G393), .b(G396), .O(n1405));
  inv1   g1333(.a(n1405), .O(n1406));
  nor2   g1334(.a(n1406), .b(n1404), .O(n1407));
  inv1   g1335(.a(n1407), .O(n1408));
  nor2   g1336(.a(n1408), .b(n1402), .O(n1409));
  inv1   g1337(.a(n1409), .O(n1410));
  nor2   g1338(.a(n1410), .b(n1400), .O(n1411));
  inv1   g1339(.a(n1411), .O(G407));
  nor2   g1340(.a(G343), .b(n595), .O(n1413));
  inv1   g1341(.a(n1413), .O(n1414));
  nor2   g1342(.a(n1414), .b(n1400), .O(n1415));
  nor2   g1343(.a(n1411), .b(n595), .O(n1416));
  inv1   g1344(.a(n1416), .O(n1417));
  nor2   g1345(.a(n1417), .b(n1415), .O(n1418));
  inv1   g1346(.a(n1418), .O(G409));
  nor2   g1347(.a(n1397), .b(n858), .O(n1420));
  nor2   g1348(.a(n1420), .b(n1401), .O(n1421));
  nor2   g1349(.a(n1421), .b(n777), .O(n1422));
  inv1   g1350(.a(n1421), .O(n1423));
  nor2   g1351(.a(n1423), .b(G396), .O(n1424));
  nor2   g1352(.a(n1424), .b(n1422), .O(n1425));
  inv1   g1353(.a(n1425), .O(n1426));
  nor2   g1354(.a(n1164), .b(n1015), .O(n1427));
  nor2   g1355(.a(n1427), .b(n1403), .O(n1428));
  inv1   g1356(.a(n1428), .O(n1429));
  nor2   g1357(.a(n1429), .b(n1097), .O(n1430));
  nor2   g1358(.a(n1428), .b(G393), .O(n1431));
  nor2   g1359(.a(n1431), .b(n1430), .O(n1432));
  inv1   g1360(.a(n1432), .O(n1433));
  nor2   g1361(.a(n1433), .b(n1426), .O(n1434));
  nor2   g1362(.a(n1432), .b(n1425), .O(n1435));
  nor2   g1363(.a(n1435), .b(n1434), .O(n1436));
  inv1   g1364(.a(n1436), .O(n1437));
  nor2   g1365(.a(n1336), .b(n1251), .O(n1438));
  nor2   g1366(.a(n1438), .b(n1399), .O(n1439));
  nor2   g1367(.a(n1439), .b(n1413), .O(n1440));
  nor2   g1368(.a(n1414), .b(G2897), .O(n1441));
  nor2   g1369(.a(n1441), .b(n1440), .O(n1442));
  nor2   g1370(.a(n1442), .b(n1437), .O(n1443));
  inv1   g1371(.a(n1442), .O(n1444));
  nor2   g1372(.a(n1444), .b(n1436), .O(n1445));
  nor2   g1373(.a(n1445), .b(n1443), .O(n1446));
  inv1   g1374(.a(n1446), .O(G405));
  nor2   g1375(.a(n1439), .b(n1436), .O(n1448));
  inv1   g1376(.a(n1439), .O(n1449));
  nor2   g1377(.a(n1449), .b(n1437), .O(n1450));
  nor2   g1378(.a(n1450), .b(n1448), .O(G402));
endmodule


