// Benchmark "c880_blif" written by ABC on Sun Mar 24 18:39:13 2019

module c880_blif  ( 
    G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat, G51gat,
    G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat, G85gat,
    G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat, G101gat,
    G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat, G138gat,
    G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat, G165gat,
    G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat, G210gat,
    G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat, G261gat,
    G267gat, G268gat,
    G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat, G421gat,
    G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat, G767gat,
    G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat, G878gat,
    G879gat, G880gat  );
  input  G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat,
    G51gat, G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat,
    G85gat, G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat,
    G101gat, G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat,
    G138gat, G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat,
    G165gat, G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat,
    G210gat, G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat,
    G261gat, G267gat, G268gat;
  output G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat,
    G421gat, G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat,
    G767gat, G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat,
    G878gat, G879gat, G880gat;
  wire n87, n88, n89, n90, n91, n93, n94, n95, n96, n99, n100, n102, n103,
    n104, n105, n106, n107, n108, n109, n111, n112, n113, n114, n115, n116,
    n118, n119, n120, n121, n123, n124, n125, n127, n129, n130, n132, n133,
    n135, n137, n138, n139, n140, n141, n142, n143, n144, n146, n147, n148,
    n149, n150, n152, n154, n155, n156, n157, n158, n159, n160, n161, n162,
    n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
    n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
    n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
    n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n242, n243, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376, n377, n378, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
    n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n522, n523, n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n542, n543,
    n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n567, n568,
    n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587, n588;
  inv1   g000(.a(G42gat), .O(n87));
  inv1   g001(.a(G29gat), .O(n88));
  inv1   g002(.a(G75gat), .O(n89));
  nor2   g003(.a(n89), .b(n88), .O(n90));
  inv1   g004(.a(n90), .O(n91));
  nor2   g005(.a(n91), .b(n87), .O(G388gat));
  inv1   g006(.a(G80gat), .O(n93));
  inv1   g007(.a(G36gat), .O(n94));
  nor2   g008(.a(n94), .b(n88), .O(n95));
  inv1   g009(.a(n95), .O(n96));
  nor2   g010(.a(n96), .b(n93), .O(G389gat));
  nor2   g011(.a(n96), .b(n87), .O(G390gat));
  inv1   g012(.a(G85gat), .O(n99));
  inv1   g013(.a(G86gat), .O(n100));
  nor2   g014(.a(n100), .b(n99), .O(G391gat));
  inv1   g015(.a(G13gat), .O(n102));
  inv1   g016(.a(G17gat), .O(n103));
  nor2   g017(.a(n103), .b(n102), .O(n104));
  inv1   g018(.a(n104), .O(n105));
  inv1   g019(.a(G1gat), .O(n106));
  inv1   g020(.a(G8gat), .O(n107));
  nor2   g021(.a(n107), .b(n106), .O(n108));
  inv1   g022(.a(n108), .O(n109));
  nor2   g023(.a(n109), .b(n105), .O(G418gat));
  inv1   g024(.a(G26gat), .O(n111));
  nor2   g025(.a(n111), .b(n106), .O(n112));
  inv1   g026(.a(n112), .O(n113));
  nor2   g027(.a(n113), .b(n105), .O(n114));
  inv1   g028(.a(n114), .O(n115));
  nor2   g029(.a(n115), .b(G390gat), .O(n116));
  inv1   g030(.a(n116), .O(G419gat));
  inv1   g031(.a(G59gat), .O(n118));
  nor2   g032(.a(n89), .b(n118), .O(n119));
  inv1   g033(.a(n119), .O(n120));
  nor2   g034(.a(n120), .b(n93), .O(n121));
  inv1   g035(.a(n121), .O(G420gat));
  nor2   g036(.a(n118), .b(n94), .O(n123));
  inv1   g037(.a(n123), .O(n124));
  nor2   g038(.a(n124), .b(n93), .O(n125));
  inv1   g039(.a(n125), .O(G421gat));
  nor2   g040(.a(n124), .b(n87), .O(n127));
  inv1   g041(.a(n127), .O(G422gat));
  inv1   g042(.a(G90gat), .O(n129));
  nor2   g043(.a(G88gat), .b(G87gat), .O(n130));
  nor2   g044(.a(n130), .b(n129), .O(G423gat));
  inv1   g045(.a(G390gat), .O(n132));
  nor2   g046(.a(n115), .b(n132), .O(n133));
  inv1   g047(.a(n133), .O(G446gat));
  inv1   g048(.a(G51gat), .O(n135));
  nor2   g049(.a(n113), .b(n135), .O(G447gat));
  inv1   g050(.a(G55gat), .O(n137));
  nor2   g051(.a(n137), .b(n102), .O(n138));
  inv1   g052(.a(n138), .O(n139));
  nor2   g053(.a(n139), .b(n109), .O(n140));
  inv1   g054(.a(n140), .O(n141));
  inv1   g055(.a(G68gat), .O(n142));
  nor2   g056(.a(n142), .b(n88), .O(n143));
  inv1   g057(.a(n143), .O(n144));
  nor2   g058(.a(n144), .b(n141), .O(G448gat));
  inv1   g059(.a(G74gat), .O(n146));
  nor2   g060(.a(n142), .b(n118), .O(n147));
  inv1   g061(.a(n147), .O(n148));
  nor2   g062(.a(n148), .b(n141), .O(n149));
  inv1   g063(.a(n149), .O(n150));
  nor2   g064(.a(n150), .b(n146), .O(G449gat));
  inv1   g065(.a(G89gat), .O(n152));
  nor2   g066(.a(n130), .b(n152), .O(G450gat));
  nor2   g067(.a(G96gat), .b(G91gat), .O(n154));
  inv1   g068(.a(G91gat), .O(n155));
  inv1   g069(.a(G96gat), .O(n156));
  nor2   g070(.a(n156), .b(n155), .O(n157));
  nor2   g071(.a(n157), .b(n154), .O(n158));
  inv1   g072(.a(n158), .O(n159));
  inv1   g073(.a(G130gat), .O(n160));
  nor2   g074(.a(G116gat), .b(G111gat), .O(n161));
  inv1   g075(.a(G111gat), .O(n162));
  inv1   g076(.a(G116gat), .O(n163));
  nor2   g077(.a(n163), .b(n162), .O(n164));
  nor2   g078(.a(n164), .b(n161), .O(n165));
  inv1   g079(.a(n165), .O(n166));
  nor2   g080(.a(n166), .b(n160), .O(n167));
  nor2   g081(.a(n165), .b(G130gat), .O(n168));
  nor2   g082(.a(n168), .b(n167), .O(n169));
  nor2   g083(.a(n169), .b(n159), .O(n170));
  inv1   g084(.a(n169), .O(n171));
  nor2   g085(.a(n171), .b(n158), .O(n172));
  nor2   g086(.a(n172), .b(n170), .O(n173));
  inv1   g087(.a(n173), .O(n174));
  inv1   g088(.a(G135gat), .O(n175));
  nor2   g089(.a(G126gat), .b(G121gat), .O(n176));
  inv1   g090(.a(G121gat), .O(n177));
  inv1   g091(.a(G126gat), .O(n178));
  nor2   g092(.a(n178), .b(n177), .O(n179));
  nor2   g093(.a(n179), .b(n176), .O(n180));
  inv1   g094(.a(n180), .O(n181));
  nor2   g095(.a(n181), .b(n175), .O(n182));
  nor2   g096(.a(n180), .b(G135gat), .O(n183));
  nor2   g097(.a(n183), .b(n182), .O(n184));
  inv1   g098(.a(n184), .O(n185));
  inv1   g099(.a(G101gat), .O(n186));
  nor2   g100(.a(G106gat), .b(n186), .O(n187));
  inv1   g101(.a(G106gat), .O(n188));
  nor2   g102(.a(n188), .b(G101gat), .O(n189));
  nor2   g103(.a(n189), .b(n187), .O(n190));
  nor2   g104(.a(n190), .b(n185), .O(n191));
  inv1   g105(.a(n190), .O(n192));
  nor2   g106(.a(n192), .b(n184), .O(n193));
  nor2   g107(.a(n193), .b(n191), .O(n194));
  inv1   g108(.a(n194), .O(n195));
  nor2   g109(.a(n195), .b(n174), .O(n196));
  nor2   g110(.a(n194), .b(n173), .O(n197));
  nor2   g111(.a(n197), .b(n196), .O(n198));
  inv1   g112(.a(n198), .O(G767gat));
  nor2   g113(.a(G165gat), .b(G159gat), .O(n200));
  inv1   g114(.a(G159gat), .O(n201));
  inv1   g115(.a(G165gat), .O(n202));
  nor2   g116(.a(n202), .b(n201), .O(n203));
  nor2   g117(.a(n203), .b(n200), .O(n204));
  inv1   g118(.a(n204), .O(n205));
  nor2   g119(.a(G189gat), .b(G183gat), .O(n206));
  inv1   g120(.a(G183gat), .O(n207));
  inv1   g121(.a(G189gat), .O(n208));
  nor2   g122(.a(n208), .b(n207), .O(n209));
  nor2   g123(.a(n209), .b(n206), .O(n210));
  inv1   g124(.a(n210), .O(n211));
  nor2   g125(.a(n211), .b(n160), .O(n212));
  nor2   g126(.a(n210), .b(G130gat), .O(n213));
  nor2   g127(.a(n213), .b(n212), .O(n214));
  nor2   g128(.a(n214), .b(n205), .O(n215));
  inv1   g129(.a(n214), .O(n216));
  nor2   g130(.a(n216), .b(n204), .O(n217));
  nor2   g131(.a(n217), .b(n215), .O(n218));
  inv1   g132(.a(n218), .O(n219));
  inv1   g133(.a(G207gat), .O(n220));
  nor2   g134(.a(G201gat), .b(G195gat), .O(n221));
  inv1   g135(.a(G195gat), .O(n222));
  inv1   g136(.a(G201gat), .O(n223));
  nor2   g137(.a(n223), .b(n222), .O(n224));
  nor2   g138(.a(n224), .b(n221), .O(n225));
  inv1   g139(.a(n225), .O(n226));
  nor2   g140(.a(n226), .b(n220), .O(n227));
  nor2   g141(.a(n225), .b(G207gat), .O(n228));
  nor2   g142(.a(n228), .b(n227), .O(n229));
  inv1   g143(.a(n229), .O(n230));
  inv1   g144(.a(G171gat), .O(n231));
  nor2   g145(.a(G177gat), .b(n231), .O(n232));
  inv1   g146(.a(G177gat), .O(n233));
  nor2   g147(.a(n233), .b(G171gat), .O(n234));
  nor2   g148(.a(n234), .b(n232), .O(n235));
  nor2   g149(.a(n235), .b(n230), .O(n236));
  inv1   g150(.a(n235), .O(n237));
  nor2   g151(.a(n237), .b(n229), .O(n238));
  nor2   g152(.a(n238), .b(n236), .O(n239));
  inv1   g153(.a(n239), .O(n240));
  nor2   g154(.a(n240), .b(n219), .O(n241));
  nor2   g155(.a(n239), .b(n218), .O(n242));
  nor2   g156(.a(n242), .b(n241), .O(n243));
  inv1   g157(.a(n243), .O(G768gat));
  inv1   g158(.a(G153gat), .O(n245));
  inv1   g159(.a(G447gat), .O(n246));
  inv1   g160(.a(G156gat), .O(n247));
  nor2   g161(.a(n247), .b(n118), .O(n248));
  nor2   g162(.a(n248), .b(n246), .O(n249));
  inv1   g163(.a(n249), .O(n250));
  nor2   g164(.a(n250), .b(n103), .O(n251));
  nor2   g165(.a(n251), .b(n106), .O(n252));
  nor2   g166(.a(n252), .b(n245), .O(n253));
  nor2   g167(.a(G42gat), .b(G17gat), .O(n254));
  inv1   g168(.a(n248), .O(n255));
  nor2   g169(.a(n87), .b(n103), .O(n256));
  nor2   g170(.a(n256), .b(n255), .O(n257));
  inv1   g171(.a(n257), .O(n258));
  nor2   g172(.a(n258), .b(n254), .O(n259));
  inv1   g173(.a(n259), .O(n260));
  nor2   g174(.a(n260), .b(n246), .O(n261));
  nor2   g175(.a(n120), .b(n87), .O(n262));
  nor2   g176(.a(n135), .b(n103), .O(n263));
  inv1   g177(.a(n263), .O(n264));
  nor2   g178(.a(n264), .b(n109), .O(n265));
  inv1   g179(.a(n265), .O(n266));
  nor2   g180(.a(n266), .b(n262), .O(n267));
  nor2   g181(.a(n267), .b(n261), .O(n268));
  nor2   g182(.a(n268), .b(n178), .O(n269));
  nor2   g183(.a(n91), .b(n93), .O(n270));
  inv1   g184(.a(n270), .O(n271));
  nor2   g185(.a(n271), .b(n246), .O(n272));
  inv1   g186(.a(n272), .O(n273));
  nor2   g187(.a(G268gat), .b(n137), .O(n274));
  inv1   g188(.a(n274), .O(n275));
  nor2   g189(.a(n275), .b(n273), .O(n276));
  nor2   g190(.a(n276), .b(n269), .O(n277));
  inv1   g191(.a(n277), .O(n278));
  nor2   g192(.a(n278), .b(n253), .O(n279));
  nor2   g193(.a(n279), .b(n223), .O(n280));
  inv1   g194(.a(G261gat), .O(n281));
  inv1   g195(.a(n279), .O(n282));
  nor2   g196(.a(n282), .b(G201gat), .O(n283));
  nor2   g197(.a(n283), .b(n281), .O(n284));
  inv1   g198(.a(n284), .O(n285));
  nor2   g199(.a(n285), .b(n280), .O(n286));
  inv1   g200(.a(G219gat), .O(n287));
  nor2   g201(.a(n283), .b(n280), .O(n288));
  nor2   g202(.a(n288), .b(G261gat), .O(n289));
  nor2   g203(.a(n289), .b(n287), .O(n290));
  inv1   g204(.a(n290), .O(n291));
  nor2   g205(.a(n291), .b(n286), .O(n292));
  inv1   g206(.a(G228gat), .O(n293));
  inv1   g207(.a(n288), .O(n294));
  nor2   g208(.a(n294), .b(n293), .O(n295));
  inv1   g209(.a(G237gat), .O(n296));
  nor2   g210(.a(n296), .b(n223), .O(n297));
  nor2   g211(.a(n297), .b(G246gat), .O(n298));
  nor2   g212(.a(n298), .b(n279), .O(n299));
  inv1   g213(.a(G73gat), .O(n300));
  inv1   g214(.a(G72gat), .O(n301));
  nor2   g215(.a(n301), .b(n87), .O(n302));
  inv1   g216(.a(n302), .O(n303));
  nor2   g217(.a(n303), .b(n300), .O(n304));
  inv1   g218(.a(n304), .O(n305));
  nor2   g219(.a(n305), .b(n150), .O(n306));
  inv1   g220(.a(n306), .O(n307));
  nor2   g221(.a(n307), .b(n223), .O(n308));
  inv1   g222(.a(G210gat), .O(n309));
  nor2   g223(.a(n309), .b(n177), .O(n310));
  inv1   g224(.a(G255gat), .O(n311));
  inv1   g225(.a(G267gat), .O(n312));
  nor2   g226(.a(n312), .b(n311), .O(n313));
  nor2   g227(.a(n313), .b(n310), .O(n314));
  inv1   g228(.a(n314), .O(n315));
  nor2   g229(.a(n315), .b(n308), .O(n316));
  inv1   g230(.a(n316), .O(n317));
  nor2   g231(.a(n317), .b(n299), .O(n318));
  inv1   g232(.a(n318), .O(n319));
  nor2   g233(.a(n319), .b(n295), .O(n320));
  inv1   g234(.a(n320), .O(n321));
  nor2   g235(.a(n321), .b(n292), .O(n322));
  inv1   g236(.a(n322), .O(G850gat));
  nor2   g237(.a(n268), .b(n162), .O(n324));
  inv1   g238(.a(G143gat), .O(n325));
  nor2   g239(.a(n252), .b(n325), .O(n326));
  nor2   g240(.a(n326), .b(n276), .O(n327));
  inv1   g241(.a(n327), .O(n328));
  nor2   g242(.a(n328), .b(n324), .O(n329));
  inv1   g243(.a(n329), .O(n330));
  nor2   g244(.a(n330), .b(G183gat), .O(n331));
  nor2   g245(.a(n329), .b(n207), .O(n332));
  nor2   g246(.a(n332), .b(n331), .O(n333));
  nor2   g247(.a(n284), .b(n280), .O(n334));
  nor2   g248(.a(n268), .b(n163), .O(n335));
  inv1   g249(.a(G146gat), .O(n336));
  nor2   g250(.a(n252), .b(n336), .O(n337));
  nor2   g251(.a(n337), .b(n276), .O(n338));
  inv1   g252(.a(n338), .O(n339));
  nor2   g253(.a(n339), .b(n335), .O(n340));
  inv1   g254(.a(n340), .O(n341));
  nor2   g255(.a(n341), .b(G189gat), .O(n342));
  nor2   g256(.a(n268), .b(n177), .O(n343));
  inv1   g257(.a(G149gat), .O(n344));
  nor2   g258(.a(n252), .b(n344), .O(n345));
  nor2   g259(.a(n345), .b(n276), .O(n346));
  inv1   g260(.a(n346), .O(n347));
  nor2   g261(.a(n347), .b(n343), .O(n348));
  inv1   g262(.a(n348), .O(n349));
  nor2   g263(.a(n349), .b(G195gat), .O(n350));
  nor2   g264(.a(n350), .b(n342), .O(n351));
  inv1   g265(.a(n351), .O(n352));
  nor2   g266(.a(n352), .b(n334), .O(n353));
  nor2   g267(.a(n340), .b(n208), .O(n354));
  nor2   g268(.a(n348), .b(n222), .O(n355));
  nor2   g269(.a(n355), .b(n354), .O(n356));
  nor2   g270(.a(n356), .b(n342), .O(n357));
  nor2   g271(.a(n357), .b(n353), .O(n358));
  inv1   g272(.a(n358), .O(n359));
  nor2   g273(.a(n359), .b(n333), .O(n360));
  inv1   g274(.a(n333), .O(n361));
  nor2   g275(.a(n358), .b(n361), .O(n362));
  nor2   g276(.a(n362), .b(n287), .O(n363));
  inv1   g277(.a(n363), .O(n364));
  nor2   g278(.a(n364), .b(n360), .O(n365));
  nor2   g279(.a(n361), .b(n293), .O(n366));
  nor2   g280(.a(n296), .b(n207), .O(n367));
  nor2   g281(.a(n367), .b(G246gat), .O(n368));
  nor2   g282(.a(n368), .b(n329), .O(n369));
  nor2   g283(.a(n307), .b(n207), .O(n370));
  nor2   g284(.a(n309), .b(n188), .O(n371));
  nor2   g285(.a(n371), .b(n370), .O(n372));
  inv1   g286(.a(n372), .O(n373));
  nor2   g287(.a(n373), .b(n369), .O(n374));
  inv1   g288(.a(n374), .O(n375));
  nor2   g289(.a(n375), .b(n366), .O(n376));
  inv1   g290(.a(n376), .O(n377));
  nor2   g291(.a(n377), .b(n365), .O(n378));
  inv1   g292(.a(n378), .O(G863gat));
  nor2   g293(.a(n354), .b(n342), .O(n380));
  nor2   g294(.a(n355), .b(n350), .O(n381));
  inv1   g295(.a(n381), .O(n382));
  nor2   g296(.a(n382), .b(n334), .O(n383));
  nor2   g297(.a(n383), .b(n355), .O(n384));
  inv1   g298(.a(n384), .O(n385));
  nor2   g299(.a(n385), .b(n380), .O(n386));
  inv1   g300(.a(n380), .O(n387));
  nor2   g301(.a(n384), .b(n387), .O(n388));
  nor2   g302(.a(n388), .b(n287), .O(n389));
  inv1   g303(.a(n389), .O(n390));
  nor2   g304(.a(n390), .b(n386), .O(n391));
  nor2   g305(.a(n387), .b(n293), .O(n392));
  nor2   g306(.a(n296), .b(n208), .O(n393));
  nor2   g307(.a(n393), .b(G246gat), .O(n394));
  nor2   g308(.a(n394), .b(n340), .O(n395));
  nor2   g309(.a(n307), .b(n208), .O(n396));
  nor2   g310(.a(n309), .b(n162), .O(n397));
  inv1   g311(.a(G259gat), .O(n398));
  nor2   g312(.a(n398), .b(n311), .O(n399));
  nor2   g313(.a(n399), .b(n397), .O(n400));
  inv1   g314(.a(n400), .O(n401));
  nor2   g315(.a(n401), .b(n396), .O(n402));
  inv1   g316(.a(n402), .O(n403));
  nor2   g317(.a(n403), .b(n395), .O(n404));
  inv1   g318(.a(n404), .O(n405));
  nor2   g319(.a(n405), .b(n392), .O(n406));
  inv1   g320(.a(n406), .O(n407));
  nor2   g321(.a(n407), .b(n391), .O(n408));
  inv1   g322(.a(n408), .O(G864gat));
  inv1   g323(.a(n334), .O(n410));
  nor2   g324(.a(n381), .b(n410), .O(n411));
  nor2   g325(.a(n383), .b(n287), .O(n412));
  inv1   g326(.a(n412), .O(n413));
  nor2   g327(.a(n413), .b(n411), .O(n414));
  nor2   g328(.a(n382), .b(n293), .O(n415));
  nor2   g329(.a(n296), .b(n222), .O(n416));
  nor2   g330(.a(n416), .b(G246gat), .O(n417));
  nor2   g331(.a(n417), .b(n348), .O(n418));
  nor2   g332(.a(n307), .b(n222), .O(n419));
  nor2   g333(.a(n309), .b(n163), .O(n420));
  inv1   g334(.a(G260gat), .O(n421));
  nor2   g335(.a(n421), .b(n311), .O(n422));
  nor2   g336(.a(n422), .b(n420), .O(n423));
  inv1   g337(.a(n423), .O(n424));
  nor2   g338(.a(n424), .b(n419), .O(n425));
  inv1   g339(.a(n425), .O(n426));
  nor2   g340(.a(n426), .b(n418), .O(n427));
  inv1   g341(.a(n427), .O(n428));
  nor2   g342(.a(n428), .b(n415), .O(n429));
  inv1   g343(.a(n429), .O(n430));
  nor2   g344(.a(n430), .b(n414), .O(n431));
  inv1   g345(.a(n431), .O(G865gat));
  nor2   g346(.a(n268), .b(n155), .O(n433));
  nor2   g347(.a(n250), .b(n137), .O(n434));
  inv1   g348(.a(n434), .O(n435));
  nor2   g349(.a(n435), .b(n325), .O(n436));
  inv1   g350(.a(G138gat), .O(n437));
  nor2   g351(.a(n437), .b(n107), .O(n438));
  nor2   g352(.a(G268gat), .b(n103), .O(n439));
  inv1   g353(.a(n439), .O(n440));
  nor2   g354(.a(n440), .b(n273), .O(n441));
  nor2   g355(.a(n441), .b(n438), .O(n442));
  inv1   g356(.a(n442), .O(n443));
  nor2   g357(.a(n443), .b(n436), .O(n444));
  inv1   g358(.a(n444), .O(n445));
  nor2   g359(.a(n445), .b(n433), .O(n446));
  nor2   g360(.a(n446), .b(n201), .O(n447));
  nor2   g361(.a(n268), .b(n188), .O(n448));
  nor2   g362(.a(n435), .b(n245), .O(n449));
  inv1   g363(.a(G152gat), .O(n450));
  nor2   g364(.a(n450), .b(n437), .O(n451));
  nor2   g365(.a(n451), .b(n441), .O(n452));
  inv1   g366(.a(n452), .O(n453));
  nor2   g367(.a(n453), .b(n449), .O(n454));
  inv1   g368(.a(n454), .O(n455));
  nor2   g369(.a(n455), .b(n448), .O(n456));
  inv1   g370(.a(n456), .O(n457));
  nor2   g371(.a(n457), .b(G177gat), .O(n458));
  nor2   g372(.a(n362), .b(n332), .O(n459));
  nor2   g373(.a(n459), .b(n458), .O(n460));
  inv1   g374(.a(n460), .O(n461));
  nor2   g375(.a(n268), .b(n156), .O(n462));
  nor2   g376(.a(n435), .b(n336), .O(n463));
  nor2   g377(.a(n437), .b(n135), .O(n464));
  nor2   g378(.a(n464), .b(n441), .O(n465));
  inv1   g379(.a(n465), .O(n466));
  nor2   g380(.a(n466), .b(n463), .O(n467));
  inv1   g381(.a(n467), .O(n468));
  nor2   g382(.a(n468), .b(n462), .O(n469));
  inv1   g383(.a(n469), .O(n470));
  nor2   g384(.a(n470), .b(G165gat), .O(n471));
  nor2   g385(.a(n268), .b(n186), .O(n472));
  nor2   g386(.a(n435), .b(n344), .O(n473));
  nor2   g387(.a(n437), .b(n103), .O(n474));
  nor2   g388(.a(n474), .b(n441), .O(n475));
  inv1   g389(.a(n475), .O(n476));
  nor2   g390(.a(n476), .b(n473), .O(n477));
  inv1   g391(.a(n477), .O(n478));
  nor2   g392(.a(n478), .b(n472), .O(n479));
  inv1   g393(.a(n479), .O(n480));
  nor2   g394(.a(n480), .b(G171gat), .O(n481));
  nor2   g395(.a(n481), .b(n471), .O(n482));
  inv1   g396(.a(n482), .O(n483));
  nor2   g397(.a(n483), .b(n461), .O(n484));
  nor2   g398(.a(n469), .b(n202), .O(n485));
  nor2   g399(.a(n479), .b(n231), .O(n486));
  nor2   g400(.a(n456), .b(n233), .O(n487));
  nor2   g401(.a(n487), .b(n486), .O(n488));
  nor2   g402(.a(n488), .b(n483), .O(n489));
  nor2   g403(.a(n489), .b(n485), .O(n490));
  inv1   g404(.a(n490), .O(n491));
  nor2   g405(.a(n491), .b(n484), .O(n492));
  inv1   g406(.a(n446), .O(n493));
  nor2   g407(.a(n493), .b(G159gat), .O(n494));
  nor2   g408(.a(n494), .b(n447), .O(n495));
  inv1   g409(.a(n495), .O(n496));
  nor2   g410(.a(n496), .b(n492), .O(n497));
  nor2   g411(.a(n497), .b(n447), .O(n498));
  inv1   g412(.a(n498), .O(G866gat));
  nor2   g413(.a(n487), .b(n458), .O(n500));
  inv1   g414(.a(n500), .O(n501));
  nor2   g415(.a(n501), .b(n459), .O(n502));
  inv1   g416(.a(n459), .O(n503));
  nor2   g417(.a(n500), .b(n503), .O(n504));
  nor2   g418(.a(n504), .b(n287), .O(n505));
  inv1   g419(.a(n505), .O(n506));
  nor2   g420(.a(n506), .b(n502), .O(n507));
  nor2   g421(.a(n501), .b(n293), .O(n508));
  nor2   g422(.a(n296), .b(n233), .O(n509));
  nor2   g423(.a(n509), .b(G246gat), .O(n510));
  nor2   g424(.a(n510), .b(n456), .O(n511));
  nor2   g425(.a(n309), .b(n186), .O(n512));
  nor2   g426(.a(n307), .b(n233), .O(n513));
  nor2   g427(.a(n513), .b(n512), .O(n514));
  inv1   g428(.a(n514), .O(n515));
  nor2   g429(.a(n515), .b(n511), .O(n516));
  inv1   g430(.a(n516), .O(n517));
  nor2   g431(.a(n517), .b(n508), .O(n518));
  inv1   g432(.a(n518), .O(n519));
  nor2   g433(.a(n519), .b(n507), .O(n520));
  inv1   g434(.a(n520), .O(G874gat));
  inv1   g435(.a(n492), .O(n522));
  nor2   g436(.a(n495), .b(n522), .O(n523));
  nor2   g437(.a(n497), .b(n287), .O(n524));
  inv1   g438(.a(n524), .O(n525));
  nor2   g439(.a(n525), .b(n523), .O(n526));
  nor2   g440(.a(n496), .b(n293), .O(n527));
  nor2   g441(.a(n296), .b(n201), .O(n528));
  nor2   g442(.a(n528), .b(G246gat), .O(n529));
  nor2   g443(.a(n529), .b(n446), .O(n530));
  nor2   g444(.a(n307), .b(n201), .O(n531));
  inv1   g445(.a(G268gat), .O(n532));
  nor2   g446(.a(n532), .b(n309), .O(n533));
  nor2   g447(.a(n533), .b(n531), .O(n534));
  inv1   g448(.a(n534), .O(n535));
  nor2   g449(.a(n535), .b(n530), .O(n536));
  inv1   g450(.a(n536), .O(n537));
  nor2   g451(.a(n537), .b(n527), .O(n538));
  inv1   g452(.a(n538), .O(n539));
  nor2   g453(.a(n539), .b(n526), .O(n540));
  inv1   g454(.a(n540), .O(G878gat));
  nor2   g455(.a(n485), .b(n471), .O(n542));
  inv1   g456(.a(n488), .O(n543));
  nor2   g457(.a(n543), .b(n460), .O(n544));
  nor2   g458(.a(n544), .b(n481), .O(n545));
  nor2   g459(.a(n545), .b(n542), .O(n546));
  inv1   g460(.a(n542), .O(n547));
  inv1   g461(.a(n545), .O(n548));
  nor2   g462(.a(n548), .b(n547), .O(n549));
  nor2   g463(.a(n549), .b(n287), .O(n550));
  inv1   g464(.a(n550), .O(n551));
  nor2   g465(.a(n551), .b(n546), .O(n552));
  nor2   g466(.a(n547), .b(n293), .O(n553));
  nor2   g467(.a(n296), .b(n202), .O(n554));
  nor2   g468(.a(n554), .b(G246gat), .O(n555));
  nor2   g469(.a(n555), .b(n469), .O(n556));
  nor2   g470(.a(n307), .b(n202), .O(n557));
  nor2   g471(.a(n309), .b(n155), .O(n558));
  nor2   g472(.a(n558), .b(n557), .O(n559));
  inv1   g473(.a(n559), .O(n560));
  nor2   g474(.a(n560), .b(n556), .O(n561));
  inv1   g475(.a(n561), .O(n562));
  nor2   g476(.a(n562), .b(n553), .O(n563));
  inv1   g477(.a(n563), .O(n564));
  nor2   g478(.a(n564), .b(n552), .O(n565));
  inv1   g479(.a(n565), .O(G879gat));
  nor2   g480(.a(n486), .b(n481), .O(n567));
  nor2   g481(.a(n487), .b(n460), .O(n568));
  inv1   g482(.a(n568), .O(n569));
  nor2   g483(.a(n569), .b(n567), .O(n570));
  inv1   g484(.a(n567), .O(n571));
  nor2   g485(.a(n568), .b(n571), .O(n572));
  nor2   g486(.a(n572), .b(n287), .O(n573));
  inv1   g487(.a(n573), .O(n574));
  nor2   g488(.a(n574), .b(n570), .O(n575));
  nor2   g489(.a(n571), .b(n293), .O(n576));
  nor2   g490(.a(n296), .b(n231), .O(n577));
  nor2   g491(.a(n577), .b(G246gat), .O(n578));
  nor2   g492(.a(n578), .b(n479), .O(n579));
  nor2   g493(.a(n307), .b(n231), .O(n580));
  nor2   g494(.a(n309), .b(n156), .O(n581));
  nor2   g495(.a(n581), .b(n580), .O(n582));
  inv1   g496(.a(n582), .O(n583));
  nor2   g497(.a(n583), .b(n579), .O(n584));
  inv1   g498(.a(n584), .O(n585));
  nor2   g499(.a(n585), .b(n576), .O(n586));
  inv1   g500(.a(n586), .O(n587));
  nor2   g501(.a(n587), .b(n575), .O(n588));
  inv1   g502(.a(n588), .O(G880gat));
endmodule


